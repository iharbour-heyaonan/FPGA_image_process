`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
R80NnScBgIZD14acGTeYZyZzlDoMDRJH97QvrM1z3/BPxjYOI5xO+RmLRE3ogivikKxeQqDB3hYo
CtT6MXJE8w==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
pzFf5UkhQCihEthT9/vXIu9qyyEco3ugn72RSG7p68vod9TXq7nS9azLrnGkzXHs3PQFBkq+3+ZG
PNN41vDN58/lK8pIjiAlp2V0xXr8ZRf/QoS3nU9pnZ3CEwxt9CGwUMks2MBnm+VSjWWRxbkUaTxZ
+kjzVWvQpUuyFFsOEs8=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
xDcafb3KrEW7vk1Eyiww/9CKbzlKF9C0uKrVBz5bHy5+6GMNsnwfCSkgxU14+VriR3jhdDN7viwB
M3a2pKPouTEOz066rknyw5X/sQ4hniBD3iUl4NQWkHTGym3kv31ZUeZYdl5ODPvzfUJOWUvkAXp/
gf4rtgV5FBbGm8qJS4jxuFSsv4rhcb7t+cae5sULvX9h7Uh0lEoAlNX3YmEW0fWj4bhIgTdzT2gk
C1ytdGU/UAnitwmujc/k+32KWV0i/o3dHRhIc31iawLLSmuBJYefDEaLG6KE8nGHeuho45Se0dhe
7kIaZp4SW1wGf7C0xxqwh1cgZ7+6eWgYBqVY1g==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OrzITnToGC+ryHZVkpDHCj6CgE4vEVrPZ7Z829783FsE2zjugDCdpipuFZ7ikbeX4Bc52TEJ4mFm
0OxylPcCXPIE74pJ186gBXkmldW4bGFMhTmUHJ94bRAsyJjr329fm+j77y2NmfbHMVOsljahWWK4
OMppytgOrZcnsnsORsbXvvikZALiCB2t+Qc4RdHc3/98o+DDvRf+gwTZNX0GMOitJmVVvqxqw6No
K3aHL26WS+5291/TUz7aF7ySSp+k84h+0omwPrcy0Xc3URWaoYbqLrWiEi22RgQYitI1tEsa+afh
tv3h9WNr+65gWTbdbwWyOz1NeXJSaNV/mc+/Lg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
riYGAyaVfIXieMgcJVFsucQ9kUNBkyzgx5CLlDibSmqSJjCaDvK63ymwoZpsGDT9Rugub8H1Y8xX
XUpLlzZGCXrlWs6NgjXfNxVpLlkmz7GswYkQ6KhUkZhRuPh0HrpJPt1ne+1pTM6fzi5LXsyTv6sn
TisWpJPdsnmBDHgM6jupb4Iv3OG7/q/NPck9K59oFLN+AyKeQ/8pEy2j7xpMiFTRlE1OTJj2mjHF
yWQWyURMafr1KK5t9Wu7YuocfKiTo0f6okHNafEo/nNpObW1D/liUJlS5GVguNNbnFjSuun9SM4T
MXhUoU0rVPqSkeCGnTpMMYK0MY5IwmbyZXn/fQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HyAIbEI1uxEAA90t6+VWFTmyUje1JDZQZoMv6A5VyFWA8tJ80b/Pwhc93aHby8xZos0WjlEANrxF
3hJ/l8XJYMVZWlVytBIRAZYGbhnMBOGo/5sjE6O2Ap0308iwfA50rb1ZITdKRqNiW+PlWkaGC+3R
QMUfNUa7cSm841V7mmc=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GUEL70ZQ78wO25wq2V+5JNZcUKzj485nYHAlIxulC+dFYZ1T3bS7X0juNGn/cdIyRbeWgA5z1viA
KyiSR064Z0BmWFsIYHfLEP1CENE6B/DkEgUM//4pBnGxH0CUe8wWHQBcyJQAxQHemECYQ5/QfTqT
96OTv0jwZ8yRjX1vKXS1qZKREGwNAsV3Kgrd9M5oaNz3PuISlyOOLoxPx9Qvu0Z0QYAzZbksLAI6
oekHTbR7CXs/P7+GCnbyf0lD6RFUyKASz8PAAvPi/+knG0A5BGQv9W8rEQ1GlCyJMbWqS7UMYIM5
Aany0Gd6zUtHqzCJMTpR0Gv6o8IS9bMCD8CICQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 125824)
`protect data_block
3YfXQv98Kli9Z1woK1QY5fYegH5TB2+PfHjJas8ZvNMVYUIX6lO1Jrxn4g63CKIL8+HfBwtE7m81
PDPpaz7nbg53aFhEprZ3xahQo/U19M+kXq20Qv369zdqX7Qj9z6BAqroBtJpcIFBebdpr6Z3RudZ
2sAnjc/crVkO432HXnwdx+g1qpR6erHM4kYzD8fduRE0rrNu46JO78EOF0pArI0UmSfFZ5pBoNbm
2CZOX6BW8yxxrosMJ2h9vhQOuLIPfAm4OwwSTe8xnQSNCnKtRPy/WxVfcWlqkeqxydu2UMdSy+gr
/N8P5fJbR5NKbX7+a5FBlPREjqqM9PsWGTLRtPaG0vVg/1EeLPOh4E8BuPY11/6K8Hyvj6S4lOHB
rafoDCNNFPgrNCs+F0b1InWk+2IPVv5vFvITYa/qFck/TOOSLn+3i6CWiTT8lufixUz6zL2JLChW
xcV0i6zBL3/6Bj/VHOV9Rl5MSVfXdtwjoILmPN5t2rxhsW0vw49VLa/Iqcm24l01VNoCslJV6JBX
He/f/BlSM5Xs66O2K7z9+JYpLeLb3MKe3PCYtO0K/a9vn+502PobfjoGXFV51jQkQnrplTtwAeH8
t7CMIkB5O0DAuvzN1oM0KIIznT0AvhD9O1ZSlQ8ayk4Me0cBWPSB7DrikyiDZ32NY1iT0zhcCoq0
MxtLf8Xk9qqPASWY4vWhe/EQNtREMxkJQK2w9SMDtXOq+oJY75VtGDFNjcQEZye9TGbCibMgRJun
Qz/tfX97XQH1qGbLI5hGB9FMi+1bw5toF0AVWlAZLnjomINJtkZlANsHZ9HTkWGUAqaTGtMNz2oE
PT0N/hXqg0pxoyhBzVDYhKQL2JeVIBGzWPKZ095dYgbKJngUPulg+e815kcN7ZVaxPkH8ObNIocW
F9mqMQ65kNrPHVTCTKfIioJjyCZK5U7R5rev+U0rxd2kvHAYB0nbd1v2dQYqD4jrzb5fm7z4F/T8
qFJvAzQVOZU3LJWF/y2Ckf0emEUZwFpONFWp7HQRrE3zfVkPMiRyZs9VlcDwjblPxyogwG9QHY8t
Ddmw5RKwdijuvCfON7hvU8W27fYj4di//Od0QHBfzWgZK3CT+0Me++rknc+xgqlHgOlxKGazbYy3
qUhn5EzlyQgalKqwQQa7Du6sWhm9eSrzvfoINWjrALsUt9kf3nKaISaLMJawd6Zh7jGMuDG5/pZj
cfwgCtwaH1Kwbl6UaPC4FKIPTtK46nuXiQ/i9GTuvnBwsyUvjTDbxBg1SC1hd3vr4+4g3aYS40ys
nx7rSia+gbwTPB++/gGTYrYsA0eWz5w7CFZYoCCJaciPK5wfTl6ulvdue74ShphUZM+X43c3X032
zW1XnplwysuO8Fv9XOCENCBYJ/BR8N21mQFS9bCBlWbBv//3C39jHAhf0zfybiKMs6Z/2S+Xq5At
Tn17SheJIIT/18YGobd4qdBRgvoUmJuVmN+vNvyxT/zKi5ue+IoOukPi1QTvro71p/R3Ql7lyLLK
wzXFy4udyf/EhPpJIXlKr1rUunvUgBcJ4ova620cZ2ryzIwGIbpT3fkWrMouAQVSPPooJi8ZeJro
HbCSbqHj/eBnQrq8yKDyEyJSt64wMyhXu7MIqpg62GfEHoilPl9NE3SGX9s74Z/Y87vcCvDpqp2D
btN+pTcSUlrFW2TNAmYw1OUP2brEgVRtlNdZF/F4wd3W2As4PHWF+XXgEigO/K35MW35+/4Gxnd4
OLlPXx+hGtLelCsEWBZLWEKxYVVS1o+t80KUn4PVrRoXvyskNjJVNFEjDb663G9h35g0qpt3pIFQ
knQWNdvebted8MDpKskKiBAQ8NYuIhULfZOQnflswhSpIPnD27x2IGi0dKTX56d9jlAtGoijGXdI
MPKzdMMdlWubEWpsWHYvK7JJVpR9UpXM4jpY+sjNm0jmbVbYXEQaXvD4U9Y9fjWWXze0IfKd1cUX
oQUP0azKPwSdJ9gOTyA6GZ/DJriMGo0u1Q/BgJCA8sirIktB6NJZDHDjM85PLgQfZ4nRkyGwXRY6
Ept1/XuTMX6pgx8Jt9SJr1TN6G8fTTL2VBGUFfzRIQnOrADYwPycty9Hnvmhg/M5eZFSFBZh62iW
BZthvlvABhAAeg74Ef6AWCIKC47KTnQ1UzuibeLDwCkDbOFryqFNPqXhlx3KBO0/9o5c4pSxuZyy
YMCpXYHLGFsHcHlOuovc60zqs9x/xGWqisvwLS5qlX/lmiLDnO+z7G7+tCl1dH+27Yw2DkYcdoGV
y3CvDzsil2qQqrH7um+DqRX1xzIJtWQlhXW8YP7I7aBkpbYKYqptXVsprGyXFuv1W31ee2XfswIN
1tB5wW1FBxaFJzg+Wt+4oJbzCZH4GmCknRcgHoGV9XyHcsXfeXY6iHlsTWEnG2/dS5r8r7MpySP+
ZIas1Jf2/MWrzqliGc9Cb8dn95RKsz42vCXwY8vWwfoeQLOAm3A+g6rMCFIjgU2o/ehbOmtDAvxA
6WA1tJX2to65Mduw+w6jtSRdanvJxsTgS05LSHiL+g6HYz8qJCzXG+naTzFPPJSK7zRuv5ODmUSX
mF44f/OvutQTKNG3kJ0JWbN1s26cbyTGtGmQNu164v2hdKpDxGvCqXznSB7OgG7LekvqMVIbrHFN
VM4HzlE2nhIMLBgoThByH3BpcZ6XkHenKDb3tyOREyU1Yame9CxfR7uxstuQHYJficsi+9mSBx29
xWESvYZAwAjhA1lZ0J260BTGVdpRuHjqxy9sbE4DWSDcTNlbIdnEBqU5GiQWmVufoWVTNvKOhoKS
dWSOcHsp6KrYYkBmqhwU9afpIUShT817iNShiPztj/IjvEgQkp6ekpFadPyNzbDNXawNVw6rAZcC
dozRm4ZNNo6w4EvvhvLEyZ8fvMAKAz5eT38c7AnpOkHMOaKl+kTe3Ogt6XqgWgMqKbzRoLf8hEWt
ootGFYo66n/Eo624676Um3Kc6flNPDC97O8MqXty1ZcjGVgjEkNnXoA6ghKtJk9weh+PE/NlhAdQ
o/M2JIFDooic/VXBznIGL3SG5RhGsgpjdDw9TVI4zQfHtQaV43OSxvy6yv+ChmyOj0XV+Cq6y56Q
EDvIjSC9vtkYRJVm1DfvQ4OcuBRPXTJUuk1ckWwmlVYZwkuHLtlhqS2Gq6GiXr+Y5MVqW08aLeXE
TIpqVfP3NaZMijl0R0JVgPEvakhSuTAV/6jdb7GwNoxJ0K0T6p1bb4aAt4EyAs8RrY4p7lDSV7OP
OAmaUjzJNUqAc6P6tyxlntQu+aam+CT0tUL9j4HggRX6z25UfIQtlw17UEJrVcEGFKRvjzOyN0A7
NjOJEtjHz+i0ZUPCPcFqxPSDOYkvttPLwgfbEF7nFzeyhBcVsmwEDaZN019ad4rJ8xniF8dyHLsz
gh3Mab2NOoT4PT1BFqIvh3n8h4VZOHrgHsrMVbiFnwB63dm1SpnXJYpj1on/UXgiGmGHfAIDgWuz
Qpk8bAKlWEcS9yKtv7qIk3B8JM6nGfSSD+3Jht2Pewb/0FOeAymNiDnU02sLOuzHJ2JmVCIiPXgS
gHZED6XmSEjjdVBbKiUJIkPZKq+s0rFb9nnwUQN+zyUJaHrGGW7kBo0vyit9mBIhHigKp32pfMO5
UwyCojOU/7HwhvJBoDPePE9YYQPP9nMQMpVrSio0+wiOFTEPEnFELR+dX5WDjR9OM7/mQyoRGyo5
pvkO5gf3dl2z9kZbWm+vQ7bBDnDdXq2dis+S4ySWNRFkEJMxGI1N3IlgoCab75EwNyOF0b+7dK2L
+Jp8LWrbQwqfA2qWJ2C9ujqfXGTAnZL0mNg+VkddPqfzq1WBMdCpuVS/78lMzwwZlNof6jD/jqBd
D6B0NnQpl1CvGMyvvNXrdo1sRh5Yx+mTgHYjCFIPF6b7appuQNw9jkzVySgqkIxUo3FOgsDpdbcC
E6zoNbDR+hRoz0jm3C4EezuoPKkwCArSPn78FcBWgV5IS/I7lE7IjzYFaRWPR/o7t6uBoM1YcFN0
KL7RYKAkQ+wm03j8TqXiVIvL+JBXnuuj34hBBFkfyfFRWnJz/wflPMQqmjYXAaenfiI6PmsBZDvr
yESAnuKtyp/vW7yWxHnKsvQCH+aqOLp9nsg1HAc0zS1nZZTOWpqJh4ubLjFNyjNJKzxJ3vYOqoUJ
Fg9CY8tmqwuNvsQmZDUqLxTsYaSB7NyumJH2Cje97cKLLAJI4Po7gVnfHvMtFArVEYlyLxPUL4U/
0zexJNRn1Jvp2cKra0QbVCSFAJbzXdzI/YqM3Ji6HcTXnWXMbJaamxxgIQVsVkTnuy9+p0q5ihWe
uGdtWfzVnszS/why9pfXEYeZEey9H50CuW2CXGt2+VRKDa2PaBtrS03CUH8i1geHG8P4B86ol9Ir
wJLyySifaXyRBoIpq0PHIWz1HhZwmAPmwkOjCZzn+lGwGdK0t69kgrJh0Z5ppr+k8WJYEa7u+8NW
bNO++ZwKxMXZHtduzTjBCabtANeFOLNEvH83oYEHkd15f95kSDVFOsg0FnyhFN6eOaXejfJk6jdA
IW9Kg7Yt/sa4yUVVYLpd5bWWmzt8d7XA3wvYBZdkGamprhKTUxPITFEMwEIiRu6OwCSQhqiMafSg
2CpAZuKRG+NwgslhbtzNMjByru6Ep1/PlPL+Y6M1zI6NkPP4R+8YwwSvNRiO9Q3r5jj8l32QSjAj
V3/IyQ3RfH9rRLv8cDQqQX2VZ8+XyShs9zkCeU7Ua57GfqD3PyWUaJkAOFhh6Vme1Z01bjH4HEMM
DplPpVSRDBbGnYO5bcmWUi7T76DP4yIVSxAukKl8P3bWJyb8+cTqWImdimo4nf6mqvdk5YiLaRtG
R/DX4MYMopjU87fOt3uwlGGreJq13nNY03eKESTjg5Dvtqi/HVCi9IQPIStsvgnpLc9ShoXssIDM
bvk+YHniS9hrgs73oWNc72UJbJLIOGiLAoIqi63p/CRCXIAfM6ZT1aNZZS5AL7rxapRTj4Zg/7HH
URCni1FjnEaLrVk4Au2Osn9h7fUh1eriYyif53fKoT3xUBcWs8QJJyLPY87FUCU8HaHQtybnbOCB
ATIl6LladFFUADd4p2MEXyxWRRoObcj+jx9o9Fjn5t5F1J+FrkseloPW1u3VF4waa5G50kN29JTV
SljG7INlIoyYRpZ6NeDi66jp3k9FpN8GyiNYbFaTh7haMK0BQ+3vRo8e/2bP3VyiK7c2uF56wpep
2BA0F4tdqmP+WPJzUMyBYa2QCaFb5CeAW9+0fsIYcGJ1G6Nw284calZNqEV8xhry09L0D9cQBsub
wmoPH3lmllZPf++DVCKAhg6uPwS7zEAqDBtZJl2KvF8YluTxoaAvD5AQ1dE0NXU5uRKVGDLgd1j1
1MsOVAd0aM17CVYvfKV5Ey9IiCbWPVcvMheQsuE/6L8q6vpKvytho/AZ3CV2RD9gTXROIuyYkVcs
sp1/zOkdIFQZryWy86xbYrNiG7z4j4lxJ9kB6R8iEbGqnG0SnAbXYLnWdm+DDxNqBXA5vn0kKQSg
sya0DpY3trW03uECmAUmUwk/NYkD4q6zQEhKpwKrf906hXTcl180P2zDukMdw2ONUrujkfRw4Tpa
6c0Bx7Yn1fQV/9I3Qar4+XQpT3epcrUaTs1dn+4YlGkmIFkAu/S9FuTp2yuRFtzJH0zRPiVas1Z6
1XoVyU+xUyI4ZTbIHWm6nFjZwv1LY8AvHtEh2N86Jo19t9ROlvGietQnM50adFPa1yi7O4fjikJj
R3vMjSd03Koq3882cEZ6/YulqPd0jTpJpdsQd7tJjkL88Xlu3fVbKJ46b7Tqjlr3ZriB3CnWZKc2
jmSWB8E6H+c14/mVFFkM5GAx0mn3G8JsZ97a2p7GYkyMsjAa8LdVrfxhqY5TOXO2msgqRxIuvIlo
kvWDexTu1nockxMW/SM7FNZHcQNndcm3g0hQj/sFmTQzGe+hvJ3wF2CJDIaldk3qZjz3Psb+cTgZ
B+GqBiOMX/lZ8mB/TWEvAX1V6bnl9zpGwYKqHkUTu9KVnnEOdc6DMPdApBoPgr5CTod7UzLykYpS
1xYAs3qsARA8L3GZZ8GLRz9jl2yV8LibC2CitXhaAcxaSFn+YtyMRse+Gz0R/RP4+yEWsdv+aCum
BPgkuOX24VQQoF1At8zNsIdR/FFounuAr6vhWu+MWUm0hcS7uAZKvzXwpBF9lNzP5qAZZe/ky5fo
Ip6WAFWo8mLksEoKUDskvaxCDQOn5eIQyf+d/Ixi4QWhUgPSlBAmeHoVXJAOYoNVmLpbDHgvU5f3
0j564H9Ett8WsAmNaLXAN0NCEE8ZaUKZfHjrt9yuNXouQqplm7qoDKIiYju+k58Xwqx0zFeNGJI4
YCYxhfuqNMWfVYXdT5tucYSKXapFBFMYkNSYk8gqij0p5mC3fdSQejBm985osEhaIs9jNGtjmJWh
6Qeg7qLz6tKh+0RArx5oTD2uRRZCP+UjeZhAerwXWPD/IAZGP2KTRIp0hidF72+CXSoKoLSV1Z86
d07/dO2DxdY5SzwDL31ycU7RaxX9RHA1aZFuOhxeounwtUW34/cnftDoncQqEZhJDPQant5/0I8v
pc2hhqABvmzpXEIjka+OwoOJPYIyVSXycXGJRmRUsRoGVaQ6gZUy3t0K1JlMhy9zKpflxwAkWswY
nrHAPiP4gDNm3fL2FKPEzlcfccgROPP7qBFXfcym7Nt8okw6yq+1I3GzflPmBHAakA3fn+HL8NfE
nArg8OLKMwKh9rWYn49ccGEaEVZAs4vrgOd/5aXLp3bqfcNbm/5JumgCIFvymFRLZu8xUigbsciv
l7XUPNREvc1bqO8SWUtVpegzfKb1ToQKjb4QI/EWWXSWfa3PgnWuer2Or/qxftm3Kobh5fylvaTF
pKxLHeF4n+vDNSjuhtTahcvBsOSzyus/oVDcBr8JMmIFuep4cqBaJN+AEc/U4XZhIfEACjWcrJKJ
rtAFdNxjOIK10hgteexNsRQCD7jmB4C8q9wnA4KoIZkJ6prBHrqjluC4ldoeQNMzsGjlEHjnokRC
jAJQiErSP6feKYojI2f4RyGkRl3cH+LPdcCY0H4Gjl0LpAAwNjT3cgS+uJLXCjWjPQFbpO9dd+yj
lUwR5vN8ZGm57V2iyQCHTIBguaub6lhupKqYTKhC6XK2pJ6zJz2QPOvm2SaQ0ID5y/3cmzDO4yT1
xlmh7EYRs3MxsnUn1eQzXt+99Py2OCTDulausUndXwzg0RaLwkZPDyI6+NR4v85gdf/6qnkilEPW
JyQGaTev+kGLYyL/IaVqWCKTrQpbUgpCyrkuz9T5FPUQjAqqaBsQDEi0ab4LYyD2zRxKTi0ENs2N
mznLzjmwFUAZxcuVJUy6cgPGiGcWrtQD+L05FN9bwg7OC0R+PUejU3Iuq6X6gCdIkyltO5b7nFeb
uNWQKbZ57JP27OKKQNGC+a5zUHNndwz2t5Xh6h2UIG6QZT92WkJJtsNTs6Ww5OscZUZVdnT9+Kzo
VxipIkEA5iCynj6c73p0XyP8QIx/XnXUJkN6eMjm92+JMJKNdOPmx/H7v1VoA0A3EoMi1vJ353g+
zn6vl6C9iXBUxLoNcisVKj/oL/nbqjJBPPIhXE7kj7H3cRGCBjK+z6e1KZq8jK1Ng1HfUnSpMVEK
3IZExPjIrQ9B5raQ279SnLZXvRo+OxdKpiRxaO6KPe9lh0lGKbexrrHf2mVx507NHFEap0lg76Wv
J6GKX2+7AkgRKbVB2ISTSU82YJKPxL0n+vAd1KsG7hTo+Z6BaAFffucPhwojb6hup9Ao0BD95mng
9VrmZypDNK7YYGzywRmon0I8Xu7HXafEg8m04Y3cHgElvEvd1O8VBrTSnebLjF3JZdOCFCs9RAC1
kzyZEhEJPUdV3GPhdZyuguyUE17eKMpduv1ghu8H5fd0k9ZBAXEmAJi1J1TDzrXcY9lqn5A8U4d6
LatM2T5MDR5UDCb0R16rnN2ajObR/SE6N4on+LnaqXuha4VNuKhMMZjSBkGVB74xOvauBJ2cmdQF
7Ms8bqI8RHHnRqScf8DP0IR9wzz1ZgRgg06W0zKeT51Jr7+lsZ8i+0RoRLY2Sk8LtlP2i81l6xzT
W/6D7KZhuclNdHavkZfGXKQo7c/4qGs4X0kBA5mM0wECwG677uqC/xK9/es2o6KoROf4hJoGyqnN
ZtFaEu2QYacJ9BqGO3lRhxX3SuRmoQPiEuL4InAZ0P8H0PcCXhkg8+mTjbm2TrLgYF/1R2zWR9+l
+54oGW+WXGmv7EGpZxI9ekEDrWrkt+C2t2saWKJNdJFaWOmU4S+fLBU3Kv/575/dfFqRp5pTygG+
/0zMjn+mGxoMlx3Gd76ajxUylIpzlbpknmhRpIoE+WPgPAoEdZpPyi4GyX33zjobwDKbRej9PlSQ
KGhZgoPLBdHWC6epKG7X/t/6PfHgSZLmYLTjy9/W+TSZqMJcLZkxVqNCbGcQYEg84ZP6TysOHury
RWO+5pePX5wG+ojzWRv0BtUckpxiQ5JObWDGm/Sa/AnsYkW1GvClYjpDfSzQ2Ji5cVoUDuzXCOPj
K5jpbU5EoT8dcXq358jUBxk+0bhJ25o7dNO5H06Z9VZ3/ggh1P9wmT3XnroyuP9PlWcF1S3uQkFj
2TnWhptkg26RUOrYUipmOgxUZFobvu93mXoqdTMm3s2f/yiTKM+nxzk9OKMw4D+nyeejyYVaBqgL
gDqc+LJ02R6xAlOcfJxu7ng5kuxEY7tIPNCf4EsC7HtJKr/PWK7R53b3gd6xsXKNsQ40rHTBOnFq
ty8+TCIuRr3FQFUZubx7EZgN5VOiQYhMwo1yZzViOqAEIaR5W+MEIdZwmZuabOt+vSsz9Y5TV7FT
DqAT7bywXqCA3jFqT1uFt5HvM9Zqc2Jjf1+fDSJauiNpo5HzLXlt1MyYp18d4Bsb97w3FQRuT+ti
hNjNWQAN22ECMotlhDdvC+xZ6NtANsINxqb0znI93amjQ+BIJIX4xUxfwGi9CFKzkOzZYA2n0pcN
OLCeYwT3pwWij2Mojq9d0ya9ihwv6A2RCiSvhcdkfQTflaDG17YXBhp9an+NHwl2uShoLKCDutgu
cD9bnIeXyQsk+j4jNyKyR9YoT/HzgCVYU5UF/UqupljoWi6nqe2ukfc4hGl3BMAocSQpk7E3wj2n
tsp0Hwll2duuRCoQwXooB6ovaHzOHZTJl2+iyEqXQoeIwcIGvPWfBGwKuOdxjS5u+bokxCfYaiDD
fRGKIp7dr1pJQyS2cHIO25ta/qoeXYUEZKz5f6uezqnAXhMQlT0J9qwI+2dxwOrIiKY2YAjLjLdr
vafTQb41fZx8mfiX6sBv7tvxaMwLhaLAh8faeJXQwDnNNdRkZQ2/5k8rR//QN3kOnC3uyG0f/cCs
8+x7e57XQ+fsqMQwNaM/+GqBj8cbxY/P1IWyzUs2XTGd6y6IL5ONBrTdJnsFFeCRMN4dYcVtMzGX
Klp+Ei/KCXlxFDMP/KUaGicqrRJbhQghvTcOCoNaDqIXi0JF/Ee6QSkCdOMeSuPkkOdUCGtabUzO
HwL9qRtTuVJEgY8zZWamn+EY4SDjMNJ7yEaaeB32ftEASOAVMaZI+5ogQ6Ng0cue8Bz+rJcoitFF
S9TtzS/h98vgncSxcBO0gcXhy7/Wufurqn+cMNgvSSN3xUCx9+glEHmcucXjv7HB0XVdC0JXKhhq
dE5vsInII6EpsPMNMZhEpI0RLQ5wzx9zLGhedynYZniePpH+3gO5lFlNfU/gXmokCEZ49hLUDdD9
okuaWSXnhmP1mcef3xNFNUZtdg/+S67mw9FEFiO6npBpXCzdA8oShHGhkh8ajxoXrKjwLXqlq9b7
pjKhFeRpBZ8BMZK08+hXBalDxa1vQ3O+XiosBr5EVlHpkWLD35qBIfL37CrpFsjfd+4d/vbOneth
c28U5DSYpB3b2CGRu1ar5zrkjJ3/kGXXY7dQ0JUa0W8gbBExeRhaqttUQUQOcy4DZfH8561TwJ1N
aBXcVPaS35dzghwDWo5U3sST9xfKCoGr4kJCZwzC4jvdmfJ22x3Vn8oPxyq07a1lECpNiCVAwT3t
2PS4T01QzU/0SdbxQGWlu2h17ntrXCKNwr6GDh/9b8J51E872/dimLPYysucIwR9w1+5Tx/vu3av
7COM+udnoDIjuEKlz5EAwigQe6wExCl1z6NYs6qJErX6C9lfoJ7yuSbEELD7ivgoKnMXcLZaV+gW
nMwcMk68w5/tSpzvDXWuJQf88JCPN7LMCwDTnxpjFev2XcVt3GMJt76t1Q0SZohccsGEltCtcC+v
Ih6SX6UMz6/JHaghGX8CSVhXc9a7r+D1sIlpfmd2XXYDunHdZF4pArinuT8oVmK7LoaWakJYY1Oo
FKUoBp5OuNcOTABwDhoGxvGWiAoBAdsolCn/E+YdLjhIy8PRe2sfg55O72AmkVnZc5ww6Mt8828x
ziM+b1URl7yrDh/ZMCM7dFbT9iqv2eeuYwLCf4Wrw8PslkE4AmKgxSjM7LHj7KPBhPXT4BjLJN4+
gcA550/Nd6Cyw1Wz7n7+SImcvxWAxvlYZs0KkRfVQgSQu6Ztiddf3OWq8WCR2lTGH1w7LvN7vB0P
JVbNSHfkkCbBNYW7kW0cNpv83QKvXnS8rWeW7xijhuBk9Xl8ePDEbzSyvABcxEzZE+fvH89l1iQE
ctluFMqrTJD4EUf1EZWE4/Bo1esXftoo0k+hpY9+fRlCq7AotIf6aua9nTmmL/AIhwK/t/MMSZgH
hG+6K0YyLyeKn586Ffa4uqMHPfKzl1Cz7J9ixFMHRFTQ2RIbpEnXD/w44k2ABqvjt4PuPehRqumb
4+DQIl4xbqkY1lqzmB/vq35lgrT1CSwIEHdc11c+oQBaM7RxdqgbV2ZipOD+BAnePIxdE9Jr12OV
2RZXAOXiODJiZkuuOuxUyMhI0GIQlHV1f1B3h8uONqyho+1FPPuYX5QAtGm3BAQrppmrxoaIqJB4
bH3SXFV8Mbb7yiIvCbyJrwg3UNQSbaydVXyt3ZpIxmUhZ27j8/uc5qoCu7ceCFDU1WHc8uYPuHkA
K3kqQWc+dSXBfoQQ1NcE4NfMg2VF0yGfUyQhC90X3hz562lNjlguTmhVuaEjdJR6vQ0LrGNjQG99
05jE+coJJ0pzuyLSuo1CUDIiED2iq7g4M8CowuJcasWSiC7hHMtYbQb+1XJ97Do2nj2Un0yUEDdW
ZGaceCIq1mCrBcMSt06tNljdxAGSfKTvOUWLIyXrJOTDXtFKOmF9hgAKoBZmJNycQCozFnUrbNVL
8zTVJTiu7G1GqgO/arzlHFbBYi6OfCVBxe5W0sPcA8N5Gw+YnxFbRQhQVz9mG8C/ilXCGqhqcVuI
UiyCWPdM7O8Qhn4MD8M57mIa0FR7fHYGNw0qim/Wj4wdyE9LWBWAQrLfDaNJVscF1aIFI74YBXr/
kCJxS1jy8AcXnyog8vFkcDgt5sGwNsJ0uBLjI7mI7DeCsMdJL5PLqiwoUtB9RNPyKyjPldYb4R0C
Hb1pRIyn3wV7+MkH1+MuPb6oJbzqki1TYX9iL5OoF4UDyUh8xXPxE9iciO77L+t5F3HfNPyJfYLI
1KZzDU3K3VOTy6K9VaQqvBNowDHNlLCSF2mgwFyrkXMmfqNvojL7oHMZ2aKmaS29mpk2dXaNZ/gY
rNd3P+zv2UTIcmgu7IAkth2a/O3mogcjCKIgazAb0Zwfx40lipT+x56KhSfHImCSycVOLPIbTjde
CKdfN4gh0v2D/AP3t8oyIeCXVB9f9mPWsY0+72dZYlljTGzNvINENm45Xn7dE6CpjtCHE5dx4DUM
JL8ZH1jqf9Apz1OC96Cyjlhp4CBU2Ef1kUG5CBGjZf8lsxTDCSVqCnqcfiqLHi6ou9NhF5IoorL7
iARzI9JPCE/l4s27eLiv055ayDLlVjDMmds+YZRRBbYZVkveVRnQBBPT4+nu9SGtFLn9yORXKfYT
OY/t6F+i1WaRzpZ0q8Y/jnGdeQNQX1DjKOyetRS/u7B7KAXCOMj+Lk9gaSOU3nhObmrtsF+KeJeQ
PUstJjryYQ+fgiDcJQ/GfqwXeXXKmABNBKlHX3aITSKXanNHNOygyYTusDVkhRUUWlfjO40JJI82
BAxFNQkCQbx+V9E4vE8ky86FZHlKwbMKZbvL5Y2ZeQyQEYzXrgES0T4He/PguQ7HYJLkipYicZ2m
3bwDN3+QZ6lbKQUUS4w2ZcTRfTt7Kz/6j5CpHG2+aGPFf47vAB+TIJy1UyIBFYCAe7rR3a11KJYo
Ql0+GE9cU483OXyX9B9Xkoz4HJCKaAaFm8R0vDJAGwmLKWJ3xUcvBwUFtcSpIsJsE7ZbWZZP5VyP
I/aQE29C2RRRJfjzNRI2tSHPHtXRGhxBZXLwaappdxhfweS/FtPNX3Wrfq7QO/RwVolkYSFa13F2
y8dSOUXsMNq3x34NBbemhIUV4H+xV7p3JgkRRvW8hUFdO3HzltRbt3R3z3vyjqmZXzCuuH1oaT/o
rH5WR+am5qOuUA3BUX1MA5GKgvDUnxBgHqWTAGfoLmI4N7fdv5RwrCgzkn3LnlWBc5lHHSYc75T2
524Z/MG9xmFiHROSlc4ufi4Q6dFxDFvEjb/io8WkBlvZtADVN8CQXcXGzZj+PAHcgJbcKSCgICLr
nqjpWFt2wgS+DYDb6ji0mQuIZnDcu3QBjFrR87Sy888NI32CTDDSFJN3MJwZew24msdRhCONFBQJ
2Y2hAiqPQdyYH3qWsSuK9MO3RqkBsKVMNmb8I4sQHuI+fHmZTJp3WHPfxtWsMBZquY8vkoCKYRwO
01WT6mivy9eubAQkPRrXdWzthA9MMWyT8KZHkVUkEptBd94lvJnSU/Jump5LSco/olbZs5aqlRN8
IHkq4R55LY7dJrNARkInehKtsRn4R6qrNqAxDNPxyKrzl/FNdp6ln7Y2XU8CWDHZxdKv39q74B1L
9QNjpgINYC1yVegZjpTzPAsaGTF2Bntye+Ta0wUBL4JEWu/sQzhh2lf838FUpTbVZJdFtePRiHye
a87Ix3eH9IDHTV6XYeo5s37ZnGYvGEr+qqMETC+aDRbDllq/IoEofzFcqhUCIN919XksLM5RMmA8
qVi8RSsdKQyw2WTuVRgOmcaSqFFtdmg14fJmTeO672jndOcZmk7iPrTxX2WXTvNA9+kl1IVwJxzk
sQn6rNbAndBoPkCRk6GfXu1Lzd40b6SfrzEOIKu0/8U1bAUyQ9h2xnaLN1BT+YNMAtDIYEn2IGSO
ho3etEn7HvNN9yXghP6MfL6OhuczCqxH9bhm1pjL34UxdKuRBLHuHffbvplB5qFxtgTVF1C8FZcB
DuMe/T983r9e8RZLZAGcVFsEgaU7XZod3+9NQeDtWdTxcpIPc/Sk3SF+dSiMfSC43eI8fYF52da6
tiEJyueH6+djR1OSAoDRgNY5LMu3njmeG6zO2+LD3NlCiqdHzmDRo6Fq0bGRRu0P3uEM1yvBO2wo
Q7OmMM5duDuHr6vBvN/9wHZjplKl9I9+Tx7K1/loi/5OZrjz0QeErWPwFRW23YlSfJHwg6w3dVQJ
S64FM/gl9S2GCx7XRrE15OQknbLtes2mzrU/1djX+sydEWx/pP06H4ZxGOwjIVvoeFu2vgK7+2gd
QxANnfTkqBVk7cpCd3/CeLElxyPJ/k5wqYaReKQDr/bQQWY2qqLDxAB47zGPBAe/PRMpx+SHL2qK
Je+r4opthxCv6Io8bsqQWMl3B81NX9108inwKqHq8H2tC8UrRqTwEB5Z5UPJ8YYhs5xCqxuhPCm8
uYX8k3hC8eEXKc4jk5iQf/E/UO6EPAQ//QkafbXIZ76cni6Jv9IicLYn4fKjn72x2IPYm6vN0E8Z
X6A9HIIzBvjHiax+p1nhYHsiMGgrkd8KxX8rls5W9PphnCbXraaQUN4V9PzyFgTAEw457hBgOgN3
RCEOuNK4CZBXlWfty30d3GnrvFGXjw0HKYZVVVDiEMale/Cr78HbhIDODpcxT6jFdJv/CWBgWBrS
zjqg8csRmaLufBHEGeud5EleHguLD0QmoH/9m3nkJs06Fxk3zRDxRlhYr8Ifo1FbwBFWQkmU4mkE
xQrO5O1CWxNL6SSPW6XzBhHbJhRG05q0WsspoIxTIDFAg7PPXKGsA8xRzySrj0hFuik5o/iVq5En
LxBL2cE7jJFD56Pa1f/E57qu4i69pLhkImvSUonk76fnzMoL5Xa176n6ZekreJ19xcykDeTWMeo5
5/0FsmmvfsWyhe9XMrwLa1iUoy6s1GKreFZFJmtu64JV8OcUROBpUHWsi0BqaQNWb8eSw0J3SFHD
zkHavogJZ2Kb/gqxv0NFQ4OfWuHIGDK0LXsJ6V6W3xcm4aCpqspH/CZso8K2caGeAYdEYDmXkf1D
xWE7FXdWhVs6EJGBxIptV5gmGWozA7CKwUa9hoFAyiuX/m9BC2mWUPNO7P7vORSuJpVZftITolrU
PyjGr4Xh3JTHi+8As9+jrX1F5PcY8dTVHSfzTMICunldFjg9eHgA9u/I6Arlm2nEMV9r/aonhMX0
PZJh6GA48ay2yFRinjGq1ru3EHPb3I67XxsnzGddSH4SHU9Nly4XYO6QOwSywH5RQNTO9ePHQrsq
E0z/QdziwxUvgBMxkm/BuF5jMG90LLpkS77mqrl+XLtR+0zjvBx3RPknn+NsOPc/Tb0TgOJljE5d
aJooFDjbKTgXD87/zaFkEIjsBwBC7v7hGJ7NvQg4E5X1OsxOrA9K5GyTzwNkrfgJ3LBF8pY5+zjq
l6nbZyb3/Jyp+HqrxmxIXgEe2p1auiv2tpOQEsFh3Z/f4bp3ULmhqrrHLa8FKxmpWbBC1UgdnSWT
nAdATrO1TCTmFfWaV2DhfzhHwJ+fXmUpEz8bpxSzA5+cXlIDOPf+74ewsUy05m5aXeE0XOpWVYn1
U9KgaY+fmuFykeUhbPw9UQJNOSab/QwtdC6g0gcxQMMz8d32XT8uSGL2BVaIhduU8GWuimeZ6bsU
WcJ53Rf2P0y056rgOTFFuI3Ozk8NT2JV/B+qsr+fEGWBhSADittSXantkVPXe5iyYOPYnaKmr57A
Y9ov4D2pd2TIWWRb9+rpZSzGHljDf0+zCzv+l/gd+729IZ3aRTpwlNuZNGd+QbKWOxOBi7pMC07f
SwPS8VCyZ/tdAr2lvluaNDqUatQ3Ggfw3e4zJVd+zRKFFppK+GAX232evyp7pEmttDNB5qod1zXi
a3BgMRClJrxIj3hMYJAe74wYEf8tnzRccnLh2hCFLUWlLgFnUtEy7msm/aiGW9FqzYk4Z3elZxVj
w8CFngwO1Wbac+ziOkCxL2aFxmkfQ1XUtj2A8aNzHBOwz+6OdFeNMMfJ2LYGYbL7GrYpq4iJoC/4
1CDR+HSCyQv5j5TQV/D9NO07tgVJVPFdhM2PVqkDAOl86FEN7JtirXuY0/ZHgdkMsBNB7CwJywDY
gnxHo1hMgCtRx6hehK0cGYMX3zFKE5wdEkR2JSa4pBB8zopBfclvN+Db8RtZGWg6q85FhSnODQw8
O14vXP3UmI2EH1oT0y7S13rimXfnTzmHIzBz9ZtdX8MT0aW/oj0LlXuRQk4YfH2zDV4i5qsuRhNF
usfpeRH3NK0rr6u4hlT+dw9JjSCklwv1EZdMfh4lNtvrrtDD/zcteAareVZ9qb8urrwqXFv/LCM5
/uZl2TmKAucK+y56ferz0rl9gpV9O7emRJz20/0+XbW7b3eULNQ9jt4zOQUX6XlGVR0DCmGBHrAV
yM+lVAn0Lj9TnARnTDTvYMRZ/a6GAkLe+GcnXBBMpYRZ1j7ETWb3c2DSfTo9QgLWG8wFJ/oJGgdP
Yff9sSXzfHWodLqXbw/NjPz0D4jFF3krSxm1E1N2ElcH0v2laj1fAVJIWAgFvsS/KmZmEkFBvsGH
sviXMu9n5PBLCZNGY9o8nvfXSBR2hKvfkPm1qPmXoj9gpDRJHTzgNlVdr1iNLcnvsdrh03Xj2Grm
wbRWsF3F2BzoEtCGNIpozLmCQJYgiXlYHJowjySCFiMq34daWwHm/9zy7SiFAJHt8D+exQSzhayC
t0m0R8sIt0MjwVL9bR/0dh+d/1GGYur6YOx5wYJzsn/Zq85c+MGCWdWpX3YJ8ksLLjej4MuiLgi3
PJ2e0wkAIo7OqzOCbmMPDHRZAhrLVyLJ5x8MfovGH2AZoTOYi+nuJwa1SEoqSA+VH+PXiIqYhhpZ
M9fN2p2n5YvIldlupiAXAnwezxFq2at7IN7HJ8Ci4xIpGq7yRZHUYpYEtFSKjqQUkz7Z3tLXDW4F
ZOsTnpB+yAHd24lenJ7HuWwEH20cpE8gAnSyFQw7njLs6oGMY9/4oWEGNm1eBVydcrSXkxsVi9Vt
6YVjxx0j8Ev0M+MwACQ7Rxs3mG8fjUi1x7Nkr7abhp8s0HPmB1AqHBLlV6aftBT3DMZncCWcflh5
OwiePr/dlWHcjfaKcYwvLYNE2O9M1HYlDFF4uHl2XLuqTfWwCVBtdhJ1Ex8yypgbwWiy8lMqQoll
umVwNUyNEN/bGmtgh/IcoJwOj2VinTQFU04h3+KgUsfWHKnz9y9iTpEJ2IOFv90i6g2ZEs7Vw+rm
Ln8EXp8PS4nkxA3YykqRhIQU8cCalEQJgVxYFpu7d4rn1vPEDyMhHCqLZ+kGfLpozZbvWD085fDi
BDsjsa63zr7taI+xfZBZPZQYvT/F2WNDGqb0jgZghhYs0ZT0AyEpdVNnBFyljsLa3HYZ3EWzZNhc
yp9zJg/8WvfxBAtgl5kzqY2buLff5j596cKVdIHh84tdw2zePHKRBAXX9MXb74JkwqMIDVQ5l32W
6il5ZuVS/1uvBVNFVVxzgmIp3QnEE8x9ECh44EAp5zGJUgF4e4n9EmEcoIoKUYVf2Aw9REVmGgk/
8bAo0v54Zuln3SwP7dkHTDjeU6F4mBaWQLw7mpBHkjH968mw5luCWu2AawSrVFWVQV3IH19mf70t
RWZocHsz5bCn5IYPYUb/hwz6meNp584v20ZaLnv9uRwYGrDtLzN0D4NNKq4j49s9Xc5dx7hm2H/w
/CcB87hfaOZl3B6OAVv4LojCe5Bm2ljcvDsgJYa8sJ7j2u3tT2/M/hlfMo/0hB3MGOaSsdaX41NA
GGTTKFofh423g7nlLCSzfKWWhkzhdIUKnepIVV8gjaasOfPzcklRDZY64HpV2IJR8oeg00US+Tg1
gppcV5KfMuiGmVFm1sLNlCPmWaw6K/lmHEq/b5XWhbrbWHhw/wJyOF+5244kM/GcpsQYvcEcqw88
qQkU8OxkMpcwGsCB8WzJaIvJoPSUC5a56HHIqgpAw/rRN7kr2ATLqL0HYXuYpML2PXHQJ6ddtbya
bpL5ulBt1PdXSWK0MAewg3We/BCL2mCYtcDtYfH8u9wGOqebe5KhFPMn3JR7W0NEaADw4o+sjQJU
qQPh2WqDL/wgLF0LjsnPB9IlDO2gtB1SRh/c1GZD3g3kkTMVWsIenlXSdcBLJzrNf1kye1S2MswV
nglvFIxtozSZ47Y8hTEeaN/MYpFlU/lpts4VWmeRoxEZ3jkFrGRJl4TmgLnc9QmfTdtytYuHelr8
0oSIH3F6g20V0AJ5IUTNaA6O3z8sHrC5rEjKI8tYFcSbiHbaY/0xit1xs4sHu25/TZKcStZcaKOs
Ledd7nAfwsfWGdvvPvHdEudts/44meGMGfxYEp4CKOLdc93PH5RteS+i0zsDARpkmIt+bgmIPaWN
eSsQf6emVRSRtwPJGuDgCIOpmyYCDMt/kNKtE7xZOibx9Gl3awnPMfe3hXGFehxmbkuZaRnjWWOY
yqi+TJkCmjHpk4nkp0KaZ3ZwGqbxqsb5JC2CzaEiOTF8knrjVTvWuiIx69ZqfsIvoMfJ6no/HPKS
fewPTZMFpC1cpTNRDEfY1eWFu/MDKP6sQ6guJ4Hu5Atra7/+AN6+c4lt0+Wj+cME7fUyvfcHmNHc
p8eovAJz+eTHLrlo8a9j1QygWPiVUg7ylqTe67wIrlSrEgIIhxljECIApeE7fEwffUAxsAWPD7UZ
uIpYWlJ4HaQYlGpNqfhOj6OtcoLq5PpyLLiE2JuqSwIpatqfxf456U1poTmJVzpmdeCHs2pCDsmz
vFsZSx2xy14TpAFWrvbaoEc64UJ+mWVTB6hTU4Prn3siErbvUqXdb8uR+rPg8EQ6LgP5mJj/UeAp
aWepR8PR5EKmzR4FjW2dZgcEW6KumNJsBJpwCfN5eC633n7spzVNHo+u9TveF7J2VR6OEdn3KzkX
LrZAbav1frrZcyvDYnTbU/FYRwV94u9pR5RQG4EoH96XADu9X9Nltnwy4TNDdG2hNJQ5FaIoB5zc
K+/b1LEh9fc1hAx4Yhp4NiWVsjE+lYqZtudOue5X5C99lMidWvFHQOM3vCguiN/Q14L4v6cdZadD
Nmdyq9yGfB1ZWEHccIVGqM4uTL6CjcRgAbaUZU9YaQ4T/jYArYUFLF5ybu28IV6Tgt/ZRpmE399m
3lG2dek6aOHw/F6TdHew5lTD/l0ml1UC6S+s7vAZ6Gj2aVGRqlA1YkpKrGwyZS1S/zlpDtH7Kblt
v+RnVU5TkxqW3zCT1S4y1dwOLU9YJc+5vtENjqh6CBvtZSr4ZNUh3Sq+Yd7ncGeTL/hZsKap47Jd
Cw4RPiF0TAJBYAxzCviz+Rhfw0xYF/U0lhZMjDAl83RzbEehN6EuRnzg95TBo/x0ISji356oH1Sg
7SwUm2uiLWrZ6TJqTC/YvCufMBXumHVrRN6un7rr7EpJEoARx4q2VVD0WzMts/BaSzQGIoeGzHbt
8VKNGOriU2KNFVlp3agssd4uiVGnonfVaF4bv/Va1mX7bybVWLdknj+fSgcFtujOsKyCf8HPyMMg
RlY2w5LFNQp8QxDEqaslXCxVF60vpglUlkq9bSEv7s0KcAfc/ja4RnskfRnTm8aYY9XXiqfjS5HT
JTiXaX8S2vZCNFYah/xlxK9yQsfYlVLJeYdCKenKwfit1tUcxVo0O89Pww6sGskB/hHd8Rkyq56W
GsSV/lNV4tFyuGkN5sfhHK8iJ1Rdcp1BtulgRVZ0dsGSktBkIQk9Y9X26JLQ2eUVJ3UofyB2R+Zj
94T0KSmet8omabU8IHZLlwofRrElz1lBPW2pD4Nh4J/JjSNq+IjvW90Ribl+mJqrk2uI3WtFK8RA
F34mIDi9QykbblITZnm9nPfHaEv7QSp3/rhVHIyRgqtsXLnK6zpLGBdz3duUqW53Tmnk4EpG/Qmh
7mAIg3o24nD/xflI6D3qylBe5cr+bWVon6CeJZTHEawZ01S0ontFojA5Xz978tMD8g4VaIzHBvIN
05XrNj2mrOYS7KgTDptxbwPhjlFgQfVLp3rG6h3eFTYRsAeINIGjyn8YnTyfxUcjdUimmNQk2JXg
ykwtLXLjq+GWDiphyD2ilkQg3aA+guw2PsSDkFS/PYlwiagA82JG2huQ+ZFmC46hezl0yC/caQYZ
+hg5vdhCtYWzJru80utAARtxHunYxEAhcaIp5+BXntjMESI8gYOpSW3M6PAn3z66nl3j38YgOUtF
6kgVNGRz1zn5nbZS9nWdic1bxW2hobz0h7Q1DGgPgUjRYDeYg6DLuIIZeuuNkwD0bnaIIGRM9+y5
nJ7yVQkmQZN3GDtZyDswZfmqKiHyFJaU4cbIlTtAchgI+JmkRdAxN9WoXwakhGGne6x61OqeaVT2
JUZG3UEqnjfp95yyeum1IhOCRBRMp+OcM15Z1hjO5AqzOCAATzW8IX8gOitEr7Ouh8gCwaImy8oF
4FhllPHu3v13lZj5PbvS3lGy2JQISuvo4xw96wsY64W4LI7Agq/QRY3orrVRAaQXeTZovRs659mt
+JTRDydDLcYKI63MPJhswj9ye6T81sQiciKBO4Nm9+YGBmJ2YSIMFSmLrLdesmqGck3kEPCeYL+4
2KOQMj0Vpd6i/8GHcZ3G1yqI7LeUM6lgOY3luBCxsLFvg+50K+rMzMtcFfeAZqqfhqjBBIpmX6xd
gVg8yiMLIhkYnXMI/4dJ3DspHp9/ZBwgRNEeTrf8mzOtLEirxd3l0VanfO1Dhz/7zvvGVQKmHeGj
jaziSHhFop5xw9RtiYIL4rulAwfXnu6kvT+DwYgtJf9MOiTRsPmEJZCSlo9WlD7zJPAAFgXXWxih
3zBPIN0EUDfL0R7+aZiWD2S0nMOWHsOpJD48Qwcfjw9qKnR/ycbfp5dRAOj+3oAPznUNPejEnOjl
IwszpDze9PZhkFGa+nAXiVwISHIzAmfZaasoVr1KlHDB9dVqgh8M4U32iGIDpj3xOU9gXUOaUoqg
d5emZgRLTCehSj6LGBpc2S9BgpF+r34w0sz7/KsPVk81D4b60FsVt5MNIrXw9oFUgGp75tIs79mi
OvxUarTs8a1QBQDoiO7a210bkPpGu8HyxnkHcnytz3XQR4MBjRUbVXgwD9pi7gy2A9qvLYAXqUnn
pPIbjl/zEYiY2fVHm84qz0B5/s0++UwJOFTLetm0BKcERX04VvAIUZqscmtsyifiZEkqISunKfQ5
7Pa3dDpPcDeEKSINwQm+14hGsqyDpcSF4SJFbXro3m22wbHCeEUDvTNICf7yLoxkvepOiQ6yW0dZ
r7RHGDz7dK+NaMyvZZbZsZO79xmj2tF9/d9QycNqe3fN5dM2p6zAoIRNGoIvvfc06NhvIuHKEQfF
vXHfMiRLock/e6YDabMB6TGHpSP4nDT+/y+jogyjz17gau1feFVIzWEWLWMEajCJ3tfSGf5qyu4y
KDbpTRZfClvZc1bfWN9ZG+QQbTC1gdOJrPAXwoz6a/UyQAu8AYUq6aNbugypoMWLd+1SN6S4+hqP
TA3bD+z7ecOHIcCVoFH+rmxvL1r3uzJX4A8gInnGLyJMXXOKSB85C8BJ3/HZz7i+19DIP3Wblt5Y
PaxZsR403bmNvUp+MwV5Io/kztPbZYYiFIAjFvNu9rSMfcdPttIT48yI8FemkiYb6b+Vem5Ss+pU
+QRCyL10PQ0YRKWSp4mKMG7HnxenNeSFZqTjtBy3DhTFasZy8XCEulZrWicZxr26HMD3t0jJlOqw
TDBnrdrislvndhQUltnFmN/aLo8+czVnvBXQYdcGJEWIrslcezg+BEMGSMdMPm6E7I7MqxNpv1W2
hS6iz1r3Q+/tfKNdmruaOSHU1DNjeYszcqTL4YAqn8FNPUdQeF6SuRRYSoVw8i7WBhh3RRHok9jz
f3NnoHGDOedY9HCfTPrb0CFZ7qfHhUMlKlbgVIsY70nKDfvMq86SMElpvPxp99H4NSxpWaTuIjgG
VCpLpjcWyRY5zhSwF0AicB+5L+vf8JwK8xvk4Rno+DQLBUsHC2Nt026EGD3rk4JQR/Ij5VvNu468
tx0aJtq8ATI0fjrthtvSFg61ctWngUNQ1NdNAw7dwHJn9TIxYG3KCFsfxIoWaLZcG20oDikk11tN
4Az2I8IzmQ2fsZOt8QaXgoPXDyvC7lLr4rsoAfNifOEk2oRI5vTmnJixqgjYk12/3LkMWiqUDP2w
n2XNPpVi+d+QmCsoETqjrpWToOFhQpGMDEy303Bo/8bxy5YhpMyu9AgZcywNmXH3DGkRi8lGx1kF
p1WpSTBbR1EJyujPXNnWjWyCjfiM7YzKXMiGSIJt8p5oFDwCvKhZWtXSR9jUI7rtnUTfrPFRbOn9
X52fFj/1Iomwr6Q+ZGKvDeBX2SwMCXsMHiHx9SgsPpOIgeWKDZ0jW2NMkpObm8TgrBKIe0q26aOZ
HDEX/ErMUBL2WRNnoSvmsyw/DIzAHThPX+THW2IydCnlUZUhdEiAEfTAfUjlZdb7ZLFMsp6HacSc
/R48dvK+CvnOLTWb9o3aSKwWRHhXQedZy6c+2YyMfhWNdYmPS2KPDJVmaKBuAhFp73jWybNIW6LQ
6262edzoYlrslQxux4E4ieskrXOjKd3ICllAY3l2FetBsN1i8okwvm4hBCAIHINn+ybcdHmc6g0R
/ufq72rHDZMpCulsQxtXlGY8fIU856C1tjMkChNrNaCYgEliZ8OkHyiBkx8ZalBlyBFO9Kn09GJ+
lklQb9vf+Y2Kp5DfnVLws641GGQupgIcE0CwtJLKTyjr5dJz1crItTK9cI78TxYDbp4uOE3cQ1+9
5L1qrTJD3sVoiXk6oJgilRPZYp6X9QteTrs/X+tW/fOFcFOYJVmWqHVquB4UFGJEvU5yBoAxqyDT
c2bPrEsaBcYBRXuk9QBA41hUbsZf9IE8u2vRUFR/tpR9mT0XgQFoewR139wCR9Al522SmOLoDajf
4LG1cIqmFbe5J1AUYt2AgMdJaglSpN6DMeBBZAUrqEFDYkIdvD+l/E4tF901V/YakS0Vg9p3NXw6
eyabV7vQmOoH5HA6CTHEkU9XwP3L5bzZxuHtbhuXG12h+QdWt+RDRTksYoytXW4OWNMV5iGBmepA
z1cwxiZ/B8iosDO5jOurEjUkxu8/+Nf/DIB2tQBWrc1HADWzN3EZtBpvevzMf7SEqLLhqPqY86U8
wlGJQGRHSDyZNZG4ThSxo9TxvfDLAGGQJEvD/82nsaRx953r8d+CeMOdWNn3JeeVN1jexhT630ft
ZHVK7NU/rpydYvL353bUrYD4G95SQ8daIf4MN7+AnDY9fyDtn3NTgcFhPnvlk5xBNAUOBosCkNlu
JfLCgGlwZFVPLZZHYpca5UCSzRPBlBUDZGc2T5N3a31BiIXyOTYuuGTMvu+QqLuqHigNgx3SKYsB
pwl7ciGLMFky25E8V8MBFUfNaS7xKzBOU3KBoQK12+g2fpofj2YtbvV3Dv0DM/0w07fCYrrjSmf0
sK3kl/LsGE/bh/oeNv6Jfr2bfzg+AB9vAXQDFC5V1HwP3ZTzBj0heL5QaQr9+K4DIotRkuP7sE8v
uF5n01TuAoXUfuBAydA5ZHVZFuqk/JjVBKijxmS5JtrhXiQ8rXHIvJtbMRBbzSGS1a1+zcm4+Uwf
DbUa6MuiAcuGP3BSDd7pRwtxYZzFXPzVtmtotHs1j6NRS/kHeSeK5iGHMp4mzvidJRwLqZ6fAJYv
avET5ysVx2C4v1KeeBoEJ82/AjHg34PTbxgwXhy+ZYFCOJCBwAYK4H2jYt22qlhi6sU/Ws/rT6/P
oC+5EUoErP5Sg78zWAzbTcLyHcaI7PK0YcbZ3x/IPOGbLd0/q6jUNzLW82kseiHFANKaWY4tY5DD
Bu3M96zEWoPm71cZq75HoeVr/on+1UVpLCcKqTERUDSoqVYDBSoXEdq/lwNYnSaoPMIQRvLUsqaV
0YSi0ICiKmtvy7WWJDBCb8SqbaSqQUJ85WJEvTMdupYKgLEvgG5tIaTWJcO32NhM5F6C3+MHUKdq
jyi/xvIQmEBq4iRzYBaw9EXguly8EKhTg5MmWvpBJfgGzK8f25E8q3oo+0BKQF13JZjO+1U9pLxs
n47b6CZxx19G0X/G/oCPPBcXc7LEaa7/hTtVaR54PHGGFJIZdJQBlck0aT9MVpgZb9RBWhc+aQh+
mX5/N0KLsKR90g6ByoyFYJ4k62/5QJqTRQPQ0vuwMupqDq6MEOAQbmz9ViW/+ftMN2ufuX3+4DQE
3TyIcncq2aa6z5JtQHW33WcKBCWporYUyHKD+A1RmPuy1QwNTzufZxPgBLipRUf2Fakbi/IUPu80
Yy2hDhSN0WCoNMUAe5VtGbld4kKcJOywHC/prC+C0l3OzYp1rWI9LTap0SwKAOLph3LAfxEyxNxS
WVyPx9qUUzMdt+4d48D8sXmIisgjBvzQWybZR27YE9KkCe+mCe0sH6OvgNiKXX3yUBElOHq+9hMu
LOh+xdcbKr//FiZWI/5BlHbfnztj1I89ItQOmmcx34rEeL3ElvkyJbhlwzcIyyswtPzgQO0kqRr/
/7mmeTsWjtlkwUqlxd9KSDhYJuoKpnX0RvV09F+f97sKp+Fp0I+bUQ9ONCn2lhQ22NeLxc9fXHM9
nRONEGlCLwfluj2sl1PsJ6mIU62jDdD9+Fr1OXmva1+T53hEBPdykyEyKwO5F+udAMghk4bH39eI
oQX27NVANUV+og6uisLvvEUlWwZP58oz1AFxMJaS7ihUdQzsrvbaj/CCyodG9ippt2MU5iMmSWXh
+wjqzRCwp7NiLHGezpLTbA+u5CamiL7OLTGIRLomprNhwL3wAX25dDTpV9MDsztjVE/joTH/Oq+R
DKywL09aylKgoQRyHmRWO5n+dOhe+xn8P/xDcrpi9Ur6WTJ3LeDjuMAlax8S898kwzBWBXclbO9W
RuH1wlcY1A7tqtVaDqiOxi61Qiia0ORjXJjwRm9mprvcZoug1X6eM2mx/7EbyDktS6diVsMGbhT7
1iBxqaMEHkcy7vYIntBqlG8mtZEHqQFmpbJDF1OmyXAJH4zE0i7ZaUMFO4Ujw+ry6671Ruq9fBSJ
VKPrJToilkbdAm2smt1keqbKZNzjds/SxtIkcRdObiQEOXk0QlHanM2sChOuN+D/4rlSMgy117Tc
jGAPOtO7vZIO1fEUqWvMrFI/EcXyQfLRZgCKuUj2xe70bkQE8VZ6x9+kd++nsB8W9bkSzJW2gjn9
Yb6D+jclL3FLHh8NXjuNinsTgoYQyqFNFK2h1/RtNArCkbsQ/rWHGP4ei8I0Sfsgyw3iwLazV+Lo
yKNfu+kEHbrVt7O70Teg3VMQk1+R6kzjKrVsAVJa/6VZp7oRfVmWQJCgu99tL7FRp9C8c73+4JvZ
RTVCh4yYlycFLdEe7JWkYTvjTR20IM+BgLmdXN8rLQQs+x0J8HDadmslD68U/2bWSZ+G2p/khp1Q
UTE97e4zUfyZvOzJCkrBrQnh9qaT8Vx5Fo8lnWpjQHg/WC145izpoBmdmvbU+l/PZR9jV47oq40K
L/bL0U9iMOPgfEZ+Wzej9NHc8rVXz5Q3PlmbfbOmNVXNuFzrsK4fiCwfSRtPFw0dWXzD3+6oGMAa
YwvA+7U+ODc/RlP9s/VUEtsH8IB99ogP7hDyDNwdpaR13bUznAxcWwNkKk8LQ9MO9WuhUb/sDhz4
mvYv7pfnlESAZ2uv0uFc3CaJouOiBzZIZcE3CGLlZQL2G8X/x6f5XWcDXcK4yevDJYRu6q0lAOtW
2Ja9pVgCd519aHO3dXT6l6WL8V8YbXln73u04s1w7ck1JheAlBQeXyPLns/thpM4+0a3jh8dpjko
vyK7CKYdIbNAJ59GaKkjI2ENFR2Ub0BOB25DNJ3V6wHG6RLGcF0rdQ20qC85X04IGvrLxMoi+kwy
Z/gwozDN3TeJ9wKs9iKWHOFw+rlGzQVqeMn6W6USVCqsZFbb+rwx9WUfRUwUNO9nPVytLZZFhzX6
cOBphA2mHsAyxU3QV5zcF73f347IU5cD4DdNx2uTYlaoBNHdGLLopkpMjwMJ737iOu1IrzNkez0d
R6BhWmKIoo4sqVzlZch5TR5iIZok/sEKOgfleAVHdIbtKmSF93xf1ZhLJuaCkmSHTdapuZevRrQ9
qtwXcUn45DKp9jFOKXlH3W1H5OVGlpj9NSvwUmdtXt+tSGSnJHKe0sTOuPSkKgc4sFyKQwqs40rU
DpXLxYkMAcv/9hwAFDn2X16xHeYOzoJ7Cm2LDI7F7z37+xB+d0V1bweRKB4oQF1kkUN75aBz7Cwr
e0Mt6iF+8x7GdHbb566nTZv+KEOd+Hd9D0yCgjSlmJbxOty26TYHi/TnRomQXxhlDg94Ma81J9Ep
fmk+wrcv/lG5u5bRT64UYb5H/RMwDgWLXbNaN7t/UBXuXL6J84+2eOqs8O1XsUvzDiPCDfA05zyI
gcoPP/BONZDlWqLctqL1FqUB2sznTxE0QNYbp35X8l0B3Uxn/8reLeMxzNWjIH4w3sYCoVQVHmNX
mFZI53fbk9pom9To+/G3NeMw6tnIZf68OcOh1ZsSW24zuZVyQZyLA9AnW8melO1wQw+DE3pYikYp
3WA3sKcbc4HuWEJNMsXrSJsHUkRdXQQ/jZqRaM/gaw1y0hXdE1zoA/O+emQGtmpAUN/oSKqiW5d9
QZb2Sq7/fO8S8a1pUwUzbumBYMrwwbJkB/Dw9pfIwy4pF2pvpNEnHQHL02iso0IAEH3j6SikJh07
uCYXzKzCJOi+vidTkoRzHSfuYU4HRIHVaVS0pJlA61CBw1bJg/z+cU2yu+6oJFnRTjDYnnVdElaS
iWwst1ed1P9YC00NplnPdwWJPGS/3Pn5uUYufONf9CoSK6vvNI/h7vgIUyG+M3Z7WTL6ZRh5gy5p
02yYHXACorO2kh+XfJECcZkupKsvXkxe5mVOtYcviEZI0m2MqvHTY7x0h9vbyq00uU67GYF0PNUv
6czLyRKFFEvb9K/+FPuOTbUqPde6uUyqs05eKK6IeEbhrpo3mUXQKiGa3DjD2NiDXklWChkW+NZu
VeZgnBB7J5K1FZhgCSKklxdHDdJPLtmD5wmUJ/zQqc5nQi0bwWKTfxkv1LMVPfSVyBhQpxA7c5jR
X2WH3keZDH9EQZKIzGZwo6gqg4ew/pdWN4dq6AbPRjUzU8xrEM+kGTELK6YsGRxeeDeSIXqcWv77
P/5+XMJGv7+oJJJRNWfu5MHquCWUm2H/nMvaoOLelTbWFuJo2yxZQxv6xICJr4vXwh+3RGC1Geo4
e2dyRcsgUhQZ20adMLkrlDRoTEHpfm2measzAL6IBizIGJpoftBkXNeSszPv7Zw9RPBsFWCJqKsZ
yrDU9vju7YbooXKCVh0D3IaZEWvuUod2OvQMRgRD4ZBCYdRSSXqC7qQFCANhqHP+JO0kVTBFhk+E
7vbeZ1tEI/7yXsEdW8B6QPmO0kOBdntWX9oKensc9pXbMq1TFoxbt6uJuEUj/TA/SLAtaaoFeq2c
vPLP8nzU6MwfWKPbq+iH2C4AwHQpb5m4A/cHTdrKV7cD8FjyQ8jnCR8R4gqSsvnwaY038H3JVC3n
rgjmKeURRE3aSSOpL/XYJVxbWX8A/FTsTVtt4bXLgB1caGGSEZ68xB3DcmK+hKJ2BATvhQzBxYP1
zv1dSFuX+R8eo6dUd3I9q+37Two3nfcGPCwqTqNbaDeTLK3WP4wnWKMJUk8gLe1istTIRTh50PRQ
+VHzDP50camz7EYjKzCzhjfL4JLO7w4fMoQ023vH/VdPFCvv0IV8ZDR3wuVKR9j9jIKzKyU4NRo7
6rOYK/P0H99tq+c/jLskhK8wbotdzf4iqU+17VnBeymlXaUGLF9RYW/RrgzFNecXNxXL3MXnf3BP
T2S83oXigv13rkKhSEE31iX/syoklae2uQgOvw7pY6cSVLUO1AGFk8Wh4xFSrKFdZgviZeHvgmHt
bzbyOZW/fvXPz3WsS77evCdMQbjjwF90+yuf0HyLUTyFGGFDHZ3IUBDsFSr7N+/G/jvBDUc5aMUd
0y87MGi/O6/KEPCquDZa7AA0TWqZnwQ2vtnoLgUSPyyU1dQzgTEsLl/UBvYWgcdIwXN8Jjg6ba/P
Hfeg/WWRdW/Rfbc45KugouKGWHgEGAWB9yLZh2IeDfTOFyx71YYoVRZKNYzsIQoch6Aw6nn1zmKo
TU8c75S1yY157zgtUL5NJfcwK/NXjN14aDP7HId/sMtyIxE7y/cwrLjnbYZamas72OcFYMqbEEXA
xm66gJL+SgzmoK/Qx5Ibd4loAnBAf0XKaoqSHrx9Bpw1yB8iMqu6HN2gEMkZcQF8DW6BWyvLqSFU
h5g442IUgt8TPuGJFNtfpHdylt+sDWS7KfRnDxW1LyxsVwQ0qqa225tGnnRwg93CeV8q1iOsKbZh
8n37K8EsteNbkjEw25e4vXpzQOQyqLS+LPNQZ6tbDtHZFZlqLkItkWWrGKTqXudWVP2rZ8yP1yx5
iNVVcm8o7v7T96e5ckaJGxBUsQYtbuLWFjXpeziSe5phrU7D63dun3cTj7ejzBShu6WHVRNY8qXX
sP0ZcZ4QdIuLO2J2jvGXg3ezhBdTDiKQ7COYDDVzsYMyA16HhI7kpkQkq/k1NU+BH2mSFsGrwyxk
eOTC+fep9sdzs+bIcVGkbhE4/ZbNhzcm9r89U7ipZ4FzQaArdFiICLsrYbCf/bEPYYZj9gBkHAJz
uWFIX6bwtQT+/RbSiz6Km5XQ5MmrHghAjdWqChGNLKK/IiY0V5pTkRVXi3rgI8IWa31HOTSI6X5G
NNz+JnGx6+QYULyPgnTu6jJB0ytyrmuno+TXFuu73/WtLHYz6+08iRLWZUUVqcBanl2t3FRK06uN
xvozb6yNaN/VHwn1AkgWYacuRZZA04sXHPtgB4rJhcbhuDNqcWsMBRwcJUqMVmKJqccZzBRwXCCX
Qk+FL3jic+S5f28hHLr1m0qS2mtPvOw4NfeEthHIR/vE5jfsvT0xusSAYUMDwUAIC2z4NKxQipWV
wuLJdIguLkwhktpaNfHFUqZ6w0dcg2sDNPGR+hsiUeqhmFVwwCuDS5Qbv61PxSbKtXD35Y0zT2ZZ
AaQkF/BMwC7ywLmo2vonr+mw6h744zBrOV1zpwmd0pWCkmHWsPlg7XezIlZWIajgO7VepSn7uh1D
xPU2690wbLI5BZLEhFMEXg5cR++JeYP/CPvZGaVkh4ArS+5abYpq7bLBrnrPqQruRQYMcGxwtDik
BcKcqAuY6bWeuAeCT5TOUjk6/v9wf+hE4Sy1gztBfWH7dpMJRg91ao0/KiDHKOVhEkXAj/i08wdi
xoTMHkFGTQtvOiinALlp7J10igb4hxkzqqqxTAIlKqtkH1cM6dclBbfVogUgQ6Olp/v3E9Voa0EU
LyY9VPeh6yGziKHiU1pdINKLA6ukt4FkyZno1IqBsW00+3hXAgXSI7o1d8em+pCscahTSmAyeadg
DmdJ9RaqlcrD8iHB1nokCv2N/ZAbxCHve20OQA03e7cXmhkn+GjUnvnqvd6tFniLhMFf1fZFLZ6k
xTbWoiBSRQsANZtNHGeY08XNqYHmqL7/VC3KXZmRDtmnvyiOAmsHHFKsBEHjf+4mv5X33STLmqSL
rgkZvv35+gf/oKU7bnA/d2POET/JtNYM81YWPUUNUaR5Cn1vSst1VlEVqNcxeTC7zvGAWzgs8zYC
eCaGpnkyc0ALh+99PogMBV4dLjLzo4M3d8Bn14noerMt51E4ydaVFBv1abmWbBnveqPoB+ajphRU
KV43q2WFnfow+daLNXoQaXfO7VSvTBArrzdwk4CCHprbEjilnMOurkTDCBz/E/ir3rW5qOLQxkPn
FNq8/p49niWSKCCDCrM9CQ+RdGWZJqUOqxr7TGgnrf6M7LFn6i1E9hw0sSDllvMjSeL6hUrqYuvw
WgW+DIvPFKWaRIgjOmN75TVIaExtAhl49+l6IQw3ctjrxnTjIcT81+46YC0wSk8uEummG7WRtqMy
I8B8S2gM/1Cl34NVl6UIzuRv1N+Z7lK92c7FHz5wS21cD6uEkwUcd63IGcaUQLJjN5YsdFmIpoxP
Ob4yv2zefL+jo9R6oq7hAmUM4A2F4+ez74ggvJApqeFYlQXXHnjGKt0NV5PqjmcC7fCZXjsRzXyY
lrblIFEErqVaVjM9766cjN7cD1Fy8/ECCREo1dmRAUFxDdgYy7nFSSbBfWgEsfhyrAZ6KQyetO44
MHTNwzmq0pphmol6rpIpadzDSxJBRM49N/S67Crfq9SFtpioc5kXOSg5ZeXosmZutTddG4ljKQ+Q
jOuUuZ+qOk3zGkFay8Bjccln5iKZjiD5bN7A48TKRIErYftrNBWAjpoqKIRK09w4cNA5fk3G7os9
cg1uGQCLlJ3xzu2q1p1esJroKRgYLUGdyGqYhYIk4bQEkkqVahz/l1aobOGP7eFEjKAPSHSFT28Z
h+suE0GXXgIlsDyO2u5QvSwuN6a1sxYfdShEzzz8g9KfErq1in8VpfIO+2jzu3ltlvNCYSVn/s+C
3uBtRZXEHfWpbnVEzJRZVwk6Kn005F26EYhYgAQ3H2M9bK0cDGQF//ySaQVSR593DlruDJiiVHkQ
HdF2YrzYm1OtuOQFfNPRro7fYUw3eFbBY1L6oTcuNZnhREx2ApwFN6Ixx0+X+EVk5PBDBKMb9IkG
lezYcBmflSiDcCxDDJZOd+TlYtVi+ptIyq9p8BmWr+3F4MOJ8PYXZbaHly/BltMwsy7oJMWrxkxX
IACwzR74pR3369bjFJYpOwWUuZcTa/ctoLr4etcnTB2eVZhC7kYMb7yVxEcvn7S41dAPoJrE7EG6
j+FgMII6qdD8IwKR9i3hvrr3LADGLZXwLtYT1EAs2NXJgLINinYdl2vrclnXOfiv9BkSVXUiKgs9
BXRO473fjntT62wHIGHHLW2gO1kuHnWfpX9xSETpQZdoSw8HuYMxZ4kpActTt2z+j/CQXb2WUyWl
OfgmauuL5DNEVuy7cLBQTSTT+cuvBP1elwnbbyab9cCsGG+uFNK6k7HHByIIj+ci5reBwV+3XR7z
u9bmrrSu4luzPWTo9/BbePA5lspkxT2kToFxDrLSk+ywJcK36apkemPMpxY2fMpCql3BKVHDLyM8
ry8BxFJKorcScSR9edBbhlebhb2pqGiPvQ6xiZ584VsMvb1PPiW2jvaHGL5dPPIuXNYV2z6xP66V
faTHDe8tJuGAGQ1ms9Pt7KNANoyyDHSi7GGZWvJQpr0u14JTug7gsRzTbsR4OJd5ruSjHhqDmH2b
x/cDZS7wkhYPdEQxEO+QE7FJUUj58B53QrSErOzHXr8KD9Md0rJy3PFum6/wapJgJbt7QDwQdah4
tNPF2trxuIL9ObNhz9WnIYxprtNH+LwRLU2AWILp57RDMXx9TtDLVx0iHCAsSVl7SYL9+iZxJAJv
trDYPT+D4ZoNPzvDEOC4sTuJ6d4Y6QBwmIKCgeeJPplWvQX3aDEun/oaN8NwQBXtRpAHq/ZBW46y
tgnyKP5DS+gjXPnt15nX4kU664DjpLGfKsts7ugykWTXdDp895N4orQh704GfsHOrHg9YYFnMrB9
P9PaOLCUTyTnZBjRVgSz35pirtwQjwYVyh30fWy8WGgG0W664vZOL/uK04VcAqUJcXcy+d4idF9F
J6F1aNBqIQTNaqbXB3EyGjSLqUdaf4Kn6hW4acgEZIaisMW1rkDzMBIfaDF7PwaFW3KBf6B3JdKd
5eVI5M1vSzo+fPXD0nXLH5U85Pl9cN9AEU1qi9hLEkF9GBiXGLqXpjBwh7X1F8Qanw4lCx9UTY29
onkEKVd/SqztSGrxK/bBNgGngoCdaRTNIkzJPLcmZNXVcglz18r+isFDYhCQPgn2G+8NW0/snY6u
BMv8ZoEWcLJXOR+pPxH9a+A/Z6swnUsH1SUopU418/OPcUWPAMPokVUyXpNqMWhTr/hOP8a27TPi
mtnscTQaIgWuN/HyKNmJXL17KuM84ICg8sCKY8ApN/Y6JIL3Stx++eFGcWYGoYBVewE49LuJzjBY
7kHIiOgxWR2HaP/ot6JPC3lk2fTflJugQA9Mdcqaqk7JioNMLDcJpAuOkoZ3wCbVgYYezFP9vkT5
n2IgmAMR7uJuosKwJzw9Zja39l50/LpDKc8iTvigCWQztcj8PsbvqEvdF138JKeKZEoniBntGwYv
dZ4mnCwThABF6OpkJeVU4KUdSnrxhpyG3xnAnr3YrMhFJyk6495/5ZGnImV4Vxo14q3/Lgt6/uVO
uZL9epXTvcb5MWWMrODPXCYU1XKttLi+w9IJgE858GaMU0G05PCWsj4kML2uuezJhzLt9odfRM5M
+7iOX4yVdH4lgLGeC1h4eNStH9yKfGK5g46CXemZiQMNWZa2pbgnJa6JDkNnlDQ1kdB87F5gpkta
QJwU87A5xxWrhrUvvOw99lrJh2YqIVWnFwCq1b7i1hAU28tWC0pvvbbr1rN9Sg9Tr30sdJ/kjdO4
u6M2nExHb6xwLNITybEfUY2H/zFvPyzh8m5fx5br3u6uWA91m6Zbc7tbWB00TdOiZOMV4wPa64Hm
ar0Ekz4SyAvQ1hFQ3FcaQFvC9nDMBKuZIJi2d5KuAbosHSizk1mzhwxVZgJwzoTNIubOED8Yul2p
DFf6NGVcKU62sVzb9P2ejY6lyY/ETHwZSCInX9hpWgG1QpLDFlQd1iEa3prOStHnZ7cHsBQ+gdTj
f5AHR2b+rtAWRU5zpOywQP/QCx4BuTyACnvvKg6E2u7uTkDLFdbZZ8bSeuqN2ZKrwzRNO7NxGxwX
ExnDNJyjZ5/ZgYxpwhJeaqSx/+V6KVtOEMUsfbW8h4/NUn/B38I8Mb7rMHD6b7e6+B2OmS+hvecf
JIT9jrUJxXZotLNA6xYdSHniLwF4UdReR17vkpRNBgfh8OozDHArs92iLEi8j1Db7sZNCm5MMC3y
Y+CQuZWoDYJC/RAXCoctEpFA4/vIk6Fc6Tjj1DcykYA19ehWDMPFaJ4BOfkHg6yq4CnutkSZh9dh
Dv+u/6kROjIk5uRSU22oUxzkPXMBoAoDwj8Iw0kOvINO1ovU3ekh2xU26h+3df1mm3H/yesrR5ij
JjdeaMKupvS22X2iGLkai6y2H/c4YyrQrtUrT/hNgfFCT9noawcx0Lvez1bXB9ftjEslmSjEH5rB
JGmKPoV6WePTxyZLcaXZQabEmXdn03sGB2HoVQ97JuUY5iWP3MvLWzVjRTmmcers0RPysCpPsiHv
0TH00ZvwOroZyeW+kfezni8sQQLvfq4T3vkcbLY/OxDVurLqnaa/pZ2rCwqH3gHQrrwq5Np9hqZe
hwqVZb2wPHOuvxDQ6Yn77HDMtDBLY9pOo1x7NmtkBBWSvVG+XzyN0pMz/3i9jdxIQXRy92QJ+tf8
jy3hfyeMkWui6eUUIy5MHgvkB7oSfwHjbna2V8VYKC7FJ/eMPW4JYRJu5MabvghNvxDggIJSDOU7
bvg2hBBPbZZ9jHhMx0zIjAdrqnTJO8OZfipY3KqnpQfFwNOaV0OG7R0Iqimy2a2RlRFx+Qkzhsk7
/HDMCzOriC7xOXjWc9tqSfAGXwLlF6PbUHt0WDppcIjSXC6ILaw3bBlOvHrsW4QuozeosLU2/oUh
oB/fUqtTA8d468KCokpJaRx0g5rBKG9NoHBtGTD9ONidR+Pv/u0QlsSH0afSR69HPFOdNtLcp6nN
DYQLfZSt/4455PXt41zXdGi0PMzUupplhTCxdN7wl2DyHw863q2Q86wzdJ/SF0UeO2BIM4RNBnTN
G6HltFpMBLV2/vboyvVPlSTVU7nf45CktcMV8i3ir7b3bj8aYxcR87By6l923ZlrHdsaf7MmYkn0
tiJRhIQV+Kzz6iyEj5RVLMKjH1CJfTsrlRM5Opna9sh1IBdsOWIR/NYjXjkdzYbDVTZBnlZt7Lwv
dqN5vuueasod8+FGkMC2Rdy5CytIOlcGJdXjZXG5h6u4FVTSAx3rGFph6TQ9z+/9q/m71vv6Qcm2
ub90ur41CvPkoZwf8aas6E1BbkiG/SvWmKsEY7EZrzSonkQaOxV51RwUKjSIX3wIX3yucm9Dt1/V
kgqSJynAHhjI4Xym22kJxTo10NtbbaN+RPBoYlf0Ml10Drr7y4h+GFL7PfTI7Franx5gg/5T9uv0
jb2IkdCw5guXejSlR3hIIeORZKvzGhhKgEsle9/6vSyo2OH7eSEFVDs7iznDHA4NotgZ0CYFG+qH
xD4XvVYHTGSResOhII0+Fl7V1PWRtLPAPSxqLIVycD4INJVftjs+tMxSpT9PStc4oKNdVn3bOGUy
5AMqSB8KqHucta/s4RXk5GIOW03bA/keHXBkXcseUWZRDP/GHz7t8PaPmACb8UIeLBY/vtjqK/Wt
CK/JZuKu3TQS/qeJk8LFs1zFm/Nyr85rdp2m65JfsuonF4KxdOlT1yeO96wQiE3ZxpihR6VHRyD2
lNvE0NynK2UQYHbuHgI4k4EY6+zQ8ZWWS4zHskdQYU6SG9GtgqqaDA+aDyXj3ocuVxbkzHAQvlIl
EguN/LUky71Uy/e+yUTm1FTdr16pCm7ffdmgTd0TIhmsaMXluvQ9QwT2XRwL2R6baNizXCT3V7wF
Q6dqOIlB3f4gEiJ7Eklke/H77H2aLzG61HX+HPGGaBC9am/i7uNmC/OIx49hWudyCt/YXp8Fmasl
9OrCvRFfGNVnKiLuZSQ6NhLMpNPUQcgiTifmypauCW0CynrCom+6yMqD9NsxXl/uyYR1STI8/wuC
fyFPKVM7oECMBb8L+jOnTXtp6f4cHlZMKc8/XyVdK3W0xijV+/fbE3MSe49oryO1y8k+ko00knH6
YPKoonxdB5Vt7PRc5+78cvr+9PAUDvKHaksqusgGzRqzbhkhpgrJR8UZLcOZz3STUIzz8nhr+4PU
CZ3FvmgSvvNS1q7zGyW5vM0cfXrGWTIcdprg2UKzn8LLvWOf+xds/VX4lpSG+f+NAWeGL/nj3ROX
DBokdQJIP0lO3fuCvbZuOnu/4hswecYoaZ46lt7eH1lN1Y9xnWVoSJfdA7zJ3kCoG6+w249DcAg0
CWz7xTnucCLEFxp0TLUBX9LTy80lHGnyAJVNy/WFMcaBbodmA/TMBJZs+WFNxeAcOkOmFd+mZnNQ
LfzeQr3Y/xffjuA/XK4EiU5J3raqy29r3AFXSdVk8fhf0C7oB4vzTadpcAKW0PMQ0E292mxdQSoM
cgt5d7p3qgqASOHRsJ2TynsPx6L2uQQv4NWR0+UzFRC3K+DTGCKq/A1E+87lX1LF6dfgHamsUMeM
V6s9yweG8s2s9l6YLiKdzkHm4chAQ47bKIrRyyS34iyLPoq0oIX0kgcE42CxgRXdo2r53NbnUx1C
ZHfLYQBvTD6F8TAliYGoOJ/ARQwBnQh6pHI20kpxwqgANbs+3vatKpZQLdbZ9i84cGuIPnMldCSD
CWOPkN4MNLgdFgSE1tHes5vIW5O7geHPJJVl6vk9Ab77zlnX3C0r5qYGXVwfOM3cynFWl2RqaXPp
iWwAnQckbVfW1hzOskIK6KQOwVtWvW79kQ4AT/dSGoPNEIFZRYfcclBasf9c03IND56v40Jn1QUJ
lYbxDh8daM4FAeYkHDxm41wGw/oGu5v+baxLpIO/wQAb1MNBbw+1taHAMo89LT57dm4V1ycGyJRS
rRayShdhgjAu9n+2E6rbiqDyZa6LbbCxY9YEM8o/3l4BwQTtWLX2Kpic49XdoCVuwZgM8fiafbPg
pwidPNOG1drkoXbYKmCKIJtCWxNEHqj8aALszXmKi+cgiih7ZAFV4ZK/cQRusa7M0hTOLt05/8NY
kDbniExRjI4kX/iWrnmJqTJHHRAmfWk8u2gt1CZMEYAwRzen3bwHosCdFg4cZX4qvFiB5znA23pE
4Uio4Bvk4S7VuiMghx4y43Z5u5vcYWcE767YmKDxPd27mNqH+ogLR9xluJpFNaEHkaoFztXN3UC+
rUH9trPRidDPhhcUVVHl+gJmwYVtVcALTSeXdKIYRjkSQW1fg8D5RSzqSIvmVU7xTRHbXm/7ltPs
TJas0lyN9wdt+F/xiG8JLGkkbXM/gNkSRuKg6x2uLK7CA52j8jI5L5bR+YmQ3r5boDFOjCrybNyF
u6XgUQd6LM36ja4G75c92fARlVZMXcgVvTFEXot7QjNfKIfUIidMmsIiZf2/Fi76/+TSxuxn3cZa
33dq1j58QESzNwkBfhrbcKGZQutEhwY56efEI6wZG4oKr1/SC/xApgSsA+Qz/2KVgj+BGjiqMQFr
EcR2JrJVTr+3EDOPBHfYRxYjYQ1H0gwTcRXOLPcvCBLFNF2SuAFzAWFW5DAZnmAQunt2utHeY5xz
iKTlc5TlisVUfZosxhM4a2ScT/8CnICx3dv3cVe2tOF5D7UoqygxmRnKVU1EhIg8hr5K5f2Aam66
6hY1yfqneg97VlRvIxghcuPs62OPlIZUwrdqG2mRQ7KbLMxfJ3MjEoMA2PIP50UG138tf9SaHxiA
HNanz3kHbQusuYPxCHEtOIE0jEGS6hFor01w5MrVXEmk+x6qS0OhiYOOZGqzu9TIzL9gtRwhzxTQ
Ok9pEfcAUk321Qcjq7CQXfiYRQdP7YX4IkrXbBukVmPQBw/QhA7P3mKqX2j64tr5lbo6rz6Mo43a
CHLOKqWH6vQnRCkKQqv6sHipFUr4psN2QtkEL1/hkort7cfGJn0sGjlYUyJxywtJvKvA0KtYZ2zH
C1dMxYC+EshB6uVfg99MfjMscMnz46g3/cUhPaFw1JMVOSCDNWMTWWgVpXbsfez1ycToBlljTa35
pim1QjgPvU24t7YlZWmOZEAGd0yZsrHAe4T46PVYISulRfwwCYgxVsP8SbevCj20n80unOb4dflc
foUm90DEuxR5BAvMs8j9TNGtiE9/uuqba8bC5aXR708ETYJdumlgHCGw+093mqwBWqk9Yu1LR4cl
i6svOGtx3UYjMLvrJ6p9wQER8KX+c5zpffRElpHbQAho7Pgf8ftAHGcd25zs8o1qZJU80NY0Wuml
HlHZQs8TPgPVeVup4X/iP3TdJGAFXSDq5kdm0nmLyI0HgQJ/QGoHq5yRAvMhl1zWuWd/wNtYh23W
T4EGEwn8scYDgFjJ/+TjYwqWNN2wYfQQW4skICJw2CDNb67vjroM+TPNZ5mdyTH4PLJU3Ut/brxD
aK54HQAbyhUlN/Lk6e2AWFY/r7K9bVcGUAtI3qHLzMNhe8GO7R9bOH/vPyJhsCOvAaHECc4HyTCA
L7Ve7RSeLhqmEvmlFrgGv7aP/t1G7HRXz2BLdchQdPnNsQQaBJ4krEvZ7vGw4+lOwYWa8p9n5ouX
B5iT/4yFtX/lgQfBqqGjfC2EI5BGzYac6F63YVybDlQjhAgZFGCs9iM2vMYfkvmqwarQSkn3f7Ev
26Mv1jRY59RGE6Z84HaKdZ6HmLUCBGtKAZIOC3cR90Px0q+udTcm/87m1xO+lOLUyxMeMJXnlon7
0tDPupiAuuuv6YhGbqFYENSeTFav8EhETCrzpwqcO3cZiAaIt0l6mrYoza8BLqW7Ss4/rwKxomiQ
iQkzu9wTGsk1EzB2vSy31AnqDDQJ463hNBr6huJdF7rckL6J/yzN5754NZufQdcVoYlG3nx8/6m/
YM95jATM+54162qHxf0OjkDmpjhAft2TmbjU0VvYiDM5Tw8v764EqexveiYPCbmQjuaJPn0Bxge7
586uEPWEyAVZeMhkDp1NqUpdC5WoZH3GJHHfN6TX7qe+PV0mI0thZhVolJce/q60BDP9C4+lfJeh
xMmtrlsmO+w2dM9To9bz1mI0Qr4wFLkCWDc3TiSZKx8RBb5aZ5vN4AJ+vQ46N61DFcYqmIEZufBa
1T/7U2Ma5zpsHUugJdZH9mFmAyxunysX7Vw6NzUNneI1k9K0cgyrSvLDJJ5MuECUj/IwrIX37mxX
GN0tLRmoRm5LhQiWCHt2R20qOIBAFmlujehJYB+122nzQgA1muA2etmOPjS8j13we/0vbkxyxWGM
LW+7LMXD5ECXeWWZQ14X37BnH++aPhEvB1+WrxaYd32SMLPkREgsQhGeI0NCjFXOMk5+4yXH7h41
rPtiwYWFhUTLvjJf6w2jN2MLVpHjbHR78hHpIBIlz1WMx75TiVaUekn5nCow1nQWpgjWwvGbP9gl
ujK/Tps/3PexPOf3DKm5Jjemb1k65B+eEHgNuti/0MHun4oTTUj28tY3iLkT3SDpvwl3ITkn6U4O
y2TZSnQAk+VqC1wq8eV7QBjRUJYmemkyC0aBz7LwC6pDtXryLn3BLwFUN/lfpUVZvNR8UtBVj0Jx
6yk1AuG8b9Z+HIEXNXx8KD4c1/tF03KM0ir90HokCHbT1qdSsi+HVv0C7OeF9ADcYnECfwmfZiQp
mWh4UGkzPv+a+B/nEWZQKRJkyt9DNC7/vioTABBZBq3UsMXNTcxx6xij1pK5y0IHfFdtIPTYRWP+
arcavVCSiM1dG9SS3lSW6/s/gUfYp5Qcq9Gy50bA8yn+dh+xXnMn7o2/7nuuw4qrfI6QgMnQ2GIU
QRcJ3MijlkspWIdZjbif6gMgzfhGEIoW8N0qfX3VYg5ZkYho0/gxnyixZ5MJI2pyWtJ4WBg07dtr
kdNiIicu/1dvZ6yiGsJexkYgZZbR7+QDULB5sdp0OGOkygQVrh0Sfj3t4bsTKquCozssZOejtCHL
INxRgHQ48Ybjt8BcaK6R6oTGFjYi3mySZhXyaNumB9moMGvTxUQZ1t7/82au94NfY0JmcmMuG5/N
fKPRL33LVwI/Ck1PexnWiQz3EiSJXtb3l/smOVawwFtqPBS+G4GOx0SCGWD1bTIl1ftG4Prvk82U
84jLDDTLP/cX+pN0wUurNtu/f9cOdTWIL36OSNZNAdZD/hdJ+ZIYdejScSHWmQVoO38Uk5tNxoRs
fI3ov7hH/TElX8M9Bndg9fiCN6O7VRmX9PRmvjBgMpOi9cFSpXED1cv0ejZdyAUYl66Vt6QPgsbE
B2mWD/NnZ/keE36e+njR/elXQFj77UJ1TGPJmd44IDC0ObodEsXLQA2BH7AQQ1JuCjTDcKxW/t4r
KxgILoaKs03Ox5EhwMmZizONV/RGqsQxC0AdYqnC43C79wwvyxS8/qvI3vlnCdtDX2PA4wrEK/PN
Y43/h2T6lPbijcn8b16ATc8swOaaC/7gqwkmbdsOrOxOuIuYlsH0uecnzYtdJdvQHDBV18NKoRcF
QSpL5X/KlBwOvWjN05hANacrkFne1AI8p3m0xlB7BMbaoODrLyy41ywfx2tLxERvPiAw/7dP65sG
/0RmtYS9dBpq5RbAmS8E85uaX/vSg7uMUzX1sPKD2k1S0RNDsZYimlWiqv2KhVj33MgX5F04qiCI
rboGTRlR79H7oG6ISPJGE1dWv0vVVpkGKXvHQ/5T4PI52MvXHipX4OWcGbx+jP56R3OWdUh1IsYi
fPdE9d1rWpYQydVCLDz2zIgLj5+IbgaVyvcPA1ndsEXM/tmBKnxiW0RUaA+2gwOPG1odRb1hNGze
G99OY8PewYeScnbZXMyvZ8ciQ3CCviHfe3n0OYU9u5TZ1FylyaEEc+Fq/sN57xDSaBSnjn1CXIkh
Ay5mvEy6OlNPWbWjFsHQrFtBqhIgI7BwrXulKEYfZQdzIvv/HlfGkulW27T8fp7VtvA2MX99LgUb
KwrHl7T3eOF5CjAdjw9Bq8dQL9XqDIH1PyyKQsDYbI2eYXvPdzcPRhzyT6aXl4jeJekE9/36fJeA
xsrUf6nIK1ANT7PgbqBvUeY6sxEBht22a9gty6h/4ujwmnw4S9Rb5eni63MSbrciMb2Or1ZdyNLj
KNQ+GrLoMYr1CH0YoyzTvBzrbmp++lr73ZdQzjpVyok0Gp9WnDb6ilTjG3EDzYeqO2RbripPGJFv
fhwEOyRBtTwWcnipBt7K7wnlUszQxkBXtTr4RF+FC6+0249RMZHG5Hd8x+HL4UXSW1KxqlLI+ycC
8gVCr6ora1lu2bVxxw7c93naQzujBg06U8o58FwzEdynTKJrOfaNSX+j3YCJflVo+Kqxw4vLYRkT
GzOk3eULbcfs557el9gBUl5VllaOeDhRVVVWHwsfZcrCUh9xu4Cx23WgR+W3WAcjC76K7aQ9yTVu
+tdAtf6vBan9pMnVV17pbN7s/1QRVRfih9v7dKKT7xeGQz21xJjlSgtPIuYL2PeJ7BcBygvDbQLg
nid1ySEvPiYF1STnLVrsOgZerCFZhHjwH2oD+raKenuRId6g1IBQZHOEXmtbiBLShVO5UcrI5dsZ
vjBW2/XzFFIayJteD5Lzi/A635NwDIXTe5zQz7nNgijr9VAfA92E0R1h6ApO0fJn7xxdQGOIFa1u
X8go230bbz2Sq6gpnfid6WLC5iaxi6D8ZayKajs9cImTcCAFfEIvZSN2/bH4hHCwLATi26hZRg2K
UBNwI9ErJl6e+QvXJb0GwKTrpimiYYJZV2fccbred626rxxK1Sv+G3QcOAbz7YLenB8wdcLVpDly
B25r1EBQ9fY83RP+G8vuWCZdBTN9F5Ac/4JraI2DRaebMNfRT9Y3eSLNF4V/AaXwv1FLCjKsIOc6
EiAImWGxadHjXKCWEWrHn4H4dka4FRHBFf4wSani1TBBioB/+vhCvhwM3BTtyC8eAc6lPwlljIov
2Ueq/x6d+SvX1jHu9/2WsjpQCi//nvCO5DePX0oVY+WgXe6RbbxnO2OeQEAslGjnBEOyFfeW5Ypf
sXn4HRkGDsnvmdPI4ZEsaTXEK7BP0hfJ18f+HvbVMbNnvPfdjvL0Zymqqk30ybgO7WlJVZS/6YMJ
q4hqMWSd9H7Fx4M9+3Iym6uQdHpuW1Gy3Kgvy1OxMYn18IuTYvpeioUMAMqqxLkN9/s2zSI7W5gK
FBvNuB3kp+0xl6UWRQcLTEk7y5pYF8+ybRkqlQ6TVEymBCmYYvLBrSE0cL6SnE215SpvaD7R0fEy
705Wbjg5l9MsSTq+lOuFYnqmsrSfqmO5+GqHoT1uuxWAi/Ehaxs5SKgrqhPhANXQtePupz7ljB2+
mnwQjtlxCQ5NS5cqJZeZPo77jPkTwy4XyuYq1y3UHhIGH6Eq+PPf0b/2C87DDv6wRR4Qx07LmYSn
JUYQEVazxyCx0VNdKbwqk+DoBORdFGnwhshpmPDEh95OOQ/ctZj8tfXvU6Zd81eGdSBHqeSypQQl
WnRcmomxMesMaJIui62LgyX4l8ZGtpRIj6M9I0sNekzmnNF7TfNIg+bLvt63l8D2v4juKsO0qT/o
PTQzPpYWNK8PZOW9OXMNsZOIVnaga3Tevic0r9QujcWUQAyeREeFVbW3XNfpO+K2qP4wqFYo8Zhb
3phNuoJisZlEH0BFsCJ+aYE1wxQFvtOuGfiYGnoAMZp55sjg9O+LuNelIH2T5KwIwa51iYOeqo7Q
3XQj//pqAblZ201JaER+Lisds2EFd63AKG0XeSj2P9vFsk2tQfidT337AD/zwJiUrmCHgaN8h0w1
Dt8qS8kK+9PpRbJpWvlZI91cWs+HQQEh/+Kbi5ooXkXWAbxMexk5OXLzpkhbFRXdnCQ6vIPBeN1P
1J8dYrXWuUCuHJ6G5QA8GmZgZSNcvqvIObOH+yGgXOKC0CdSRRfOVDkJ0A9Zal9SrzI3mkJSg0bs
PT1ngKGsO3+JW7SYaLudvluiJ6t8umo8iz6MOEz4nUqruAmui8FgAthLUScXdrD5+esnfIgVjeNP
+zuI9PUHQwq/WiDPzA9Cv0ibPXT2fF2qjXGJxeccdWaqWWMl4bEEvmlTJU21J7X9opWmeOXHNxzG
RzGwraiNjIMGQT9PcRM1U6GtuYjqPp9b7ETDO0sGInQrlOkXClla8CO4MYtkSRnBIX3qtT+NkbVH
nE+cU+zkhv1l3sfzUDHTXKvEu6qNxn2BQOSWThCjNQCUTLl4ECamm80SHMRo4IkgyVDrDJdDLT5s
HCL3HrzUFG+oAWTa5WeiaB8PdaZZv0JLmSM+UYnJWK9DNIpdgUgqBg/YVUSnIz0y8YMT97KDp4oK
+rmv1wtmm2gvwpAkIiXx7Tk7VW0jomqxAVdeCF/9+t1yf/Jd/FaiO5t/paPk7Qggh9uRHfb4Xoqq
O9vxFgTDWhm8Lbg9nd9yozVnYuZf53ofOyEZVk8iccv288DUE3aejfxQ/i4H0JWXf/Kk5DJn2G9Y
RA4PjdfbsKPjpF9PsSpsYBtqayysDfSBJvxvppke91JMbMLXIooAvueqN09OiJR2lyiJT03PjaWP
YUDWTP44AmQCOqrrVxuDw55TCWUywQyw2mLMRNI8s+3ZEqU2K2O43oSdW8zlauc0/G1oFnZr8agz
TjMVKTob0PRafE+vvyQEl9b1a8euCb6h+DDqmnsYgvmzlMLd0B5nKyXJ4ZCu6tDXu+jbB2p9JXSR
hQgIK00H0zeJI1ty+XgLelCHu1XDVv6X4bO6ZXbBj0Y1gEjSae4z8c4J4cRLZ0NC2rzHWUr/SJsB
/dszMaGgM6V7aXomB6PcohoR4JBI90ilquNhONCuCFHs07lL4LWx686FLi2vGbVIoC1oTbi1tXHK
kRwRXGxeOT0nALGpoaJjO/f4W6nE9avLPsxh06VHwuzsU7ei/0EBaBoeF2lbKFPJIzBdNIbC5t6y
K7SABzWi2olrU403HHYa5pGbg3DTsymrJinToyx7Og3TjFjUpSOMQsNZLDkL83ArtzuLVYR28uE9
QXmNzj55kkR0mpH5lRnnluYJKrpWQYzJ0SMsG/lzGMkF7vAjVvGmoRMsD5HK/IDpvwFmvic0JZ8+
oDCzz/Bix6w2yzZ+J3sson+xguq2p7k+QqoaHBXix+erBaJchPegi9aO5QJeNZ6gW1RUdpPBRJ/v
Ewd0URVq0gwEzKMJDDQ0WtBUkdDc6tA6mJuN+YFlTb64SqhxQNjjOVu+GeiJNWvqsxtJ8eEIGsL3
sK6Ki3sjR6EvbDzjnq7mlCqxTdVSj3Yt2zntWs+AYhm4oRyOUX102Rf2Xq57MEhQT5THHvdtxl88
bgM1YjhnwgoGuR5yWhuG7JZtBtBOmmChXhHYjnBR7YAU9iWxvyygjl+C+25LgiRmGjgwEwb8MJlV
1B6scffJHJ0ARDedEsWpRFnppZh+jLB8V8CshwVVHIk5eUNf1G1fzc3DQtnEh53fqdwTanxbcdGP
nbYkWrMnRUEt3AzRO/g2G7GWjCCdmXm31fLqDd4I38IY6mGuPpsd576YIydB3Me9RGyMm5CUrgLk
uMkuN9zDSe/MpqevRKOf8mKiUAYO97zzFy1GRw4Hy7ZBsGrHTbCKoG6NI0LanzxWT+2r/iUdNdOR
cn4HooKYjlk2dG1q+oJ86vF+DuCMK1j6nmQo71q3RoI356iQEwG13Prn5suQrrKgAZiDXgdiIspq
nTW+tFH9Gv/XB+Q3qDLx1wDhfq23anMtfHPiBXGMR7OjTivA9yyENmYa5ndBkenTPW7/K+c25d1d
eSohHkAv/g8VthRBk+J9+x/MojvisWxRkC1nvH+K7AxES7u+qknvmcgm8vzewLYAcHluRUTDk3B+
pi11ALiOzb3M9kzdrGa8UKlTtkBZP0d93AtuLp83IkPj1tpi9nnVgxt6N/c81g1a5+M3Jz8U55QH
vQSBWp7LBYLAP1pfBQY3t8LuxaiIyjh+GbNHnLr8HUUwPyXNPQ9rwp5nIb5tAFY0RSy+rsmDTEJh
ljGCNAKt+2UEQt5zGDpDv0G0OtiJsTGXvPbFnnuUYnhjnUZmCIH6rlwGGjefVyfdZcGq0yGj0T9K
O7KQkvj9ZV/i05JgWxz5lg3b3jZOPo59xCQrRsNaOZonIKj2Wm03PuZgWIzsIYi0GPf4YaYSJFQG
JBwu71DCZGLWlRtdYTngcdEYQCfs3kq8Dtnoljieqgvu9hphunDqxew6HSqnW+lCywj6+3VAL7Xh
WDlSSKos3+rnZXOjGAl4oiRdOUrte9My3e1MmjlfnwpkQ19gHlh3jWoZONOwFN/gCK+1QZdXb78B
rQDtTjK2UFKYslppoHWOeuXw1/v4MiDNYzZYg0Q7q+sUGHk7NT5c2GyGXEyybQU7Nf70yFdSGlEm
SjjwWrip1wFXOs9pf+sA/DXN5h8Pbbmdc77UmuxZhHp9C+nRzdQ4bDqF2JBGwZZIyB4mE2b1gQN8
k9ZIoa3fkK/h0UbztUGUpTXYoEr+Ou1EiQ5jZtJ3rrvre+NAC75uv9k5gcYMypHIIhRNeMX3OkAf
1X10OER3PPHFH/MgQDTqHTAxH0WckauyE8YEdgcrUb8c6brQwNBazsEbwPkkE5YIZdOmFVjzvvO5
ZSlkQ1Hh0gZ16ZE2Fc7qt9sndGMU21VYCPBV631v1tyT6RUsfsjL4MaZM6JH8BNqkwx6QOXqVqzV
ws2HPuMIjjptco4myoyYmx/qRZ+dtOhL3FGdTpsg6sAjBQ6/D1lmNn4FB5RoDneeXpYkgZ37QHor
Eh73b/wiNGyikKc/IGKFzHG50cZGX6X6Htd+Kp6QQzgeKtuvKvnPO7Gfr4QO3BWw00hAcKc01cML
DJep3OnKz63vGCuJBeXfn7v7Rl8keDzovAKa7XcJRMv6JEPgrV4Ka0L5y95veW+vvBbjFvV8kBan
PxVEtA20CPV0IuGxgMwp4IDX8KQWgWGSrfuzchmIEWKepoe8RIPMa0gI1Z0OJIq473DKlmqnRito
MuTjaBIBo1KbILEmclVyq7j8dCRKCHDqjcOGxijJEMc9GIjp/1GiJz1aGAcFwYA6MvX3BFJ+Wvz7
ClvgENLRpeVFJ7Nq+c3a4fU+9ObA1mQEsA9psqoM0U31fzz4kMFBMbpf43wqx32T0nHItPe4QXvf
kCAO4Gb45Z/5NL1wtH7no4FvZXE29Ba5jfaaMcMqFE1QY46FobwK3jwCPnLbJ6Zm/16cdddOKIEF
CNrD+3WIrNTqyHmHJnsPGPsF0/aqh4Qyzs7RQkCHDy5wGEYGYkSS8Uv3jdHrJMWQvnOAl7rymZnS
9mIsAS7h9GJyoGDsRDJ59drAdrehqSa9fObLvvmwSUFNuBDEcWcyjkvyRGtKpvM2m4O92zQj9aNM
Ea/XtPfQw2q/G7WWJShv2eOuWzAwTud/qGj2malNJO/QoMlvUCr7OC7Mpskl9rOYD9Jeza3cZTxx
0uzvSc0Q/TcnGMMElESAznp8zbMgOk85bHb6bklSkecOgDhdxKop6A9yz9bJRNhD07r2Ow/GQ8N5
jn0JSNx993o0oIzpUv6qEFD3vN54NudF40r3Qh8HZ6YKj4U+uj6Td3K2Hdd8oFzeXpFvj9sfbJdT
adzs6RBJucrpSzDWfOOg8PYwQRHiWWxVLH/wCHdR/Q9Mf+tyndsEfPScXPUS35KU32I185We5kcI
j55wvP/uoythb+uvwrVSAGRbZP/8JQQDVrdHOg5cmItGrglNKaxHAFvJhpRHjCKGz1zytpYrSfmv
nEOFtksLfnoyMbudiONo3W7ZPOhnhP7k5pQ5EMbJO7pHtQ4za/3IuaGbjluBXQYpXcDX6NprJY+0
nuE/XkOolMSBt02KKGRwjt0/oLGVXhjK2A41tWLW9Qz4L8oRyU1PYj0b3ut3JiXl88xBRHgHYic2
y4IKiQ/shbvaUC72ANm59wsNeJ8LUi92nB//7qiykL8rasRgvaPnaUKPc0Xs21FbriLUnkqEL/y8
lND8gOsl1NYIfIpkJNu2YEG6RHjUs8haonrPHxlOcI9xj39EcdO10BueHTEhNfj1gSRDxpuFODja
U1BR8WYe8bKiaDMhTKhvpK7GLO0odX+QrqMCdohkNUU2QFtNWhILd54Sf9hIpQx9GAk3x+P48pq3
CjrEPffG5lEWISME6Z41zrcq22Fj9sZjIOlvG6C9R1jWsprtfBbOlT16Pt+bejPuvY58xY0S9ADo
mRfqOgbxmDGkdFud1NLgBptmZRrD0G3XrAYQ9AOs63IE9X5oyo3Xr70patSWFehGxwTJeWHxcs2D
27pWw0iObGZDpqRS3EeUXbcYuQUGAOJ8RyHeLm/1FVgRoyUxBk2bZgtTQPz2xrUZvVjYVSZ7DKIl
wSqoPcaYk/F9Eh796smklt9X+TxgRGmMxF3WvunlXKrfYulIvqZsO0JiFpZULydJEoOK1wfM819S
zGV6nIcmX78FyysHccGzkiuro4Y2QtbjITKop/g5KlFR9NAAiVkQZ2YjIZLzR3aeGDwsemEMds6h
NeqnmJ4mvQyJ0X9ZLOz3EEca25khdFdofMXxa6FGDSE/kOHLBrABacrrUn0f4FTqLs5HFHe5QqwZ
OKLylZKnxkHMM5iyJvIGIvgpm5pWZQylrX4PVNPVfaNSOmabDUyte1kOv9erWlyQvz8bSkOi2mF3
EFM6utUBl5Zq8cmI1Q6YGH358ZepY9MCCKcIfnJAimO19Bbu5jsCz2qbmOghDMre1P2ymcG4XA2S
buuDcmF9eHNyd0KDGXIBeJjHmRtuOoEeQL8Hxn4rld/T9GkoZtAzfqq7J/jx4X3Zgx0z7pcNHF1j
e35bHVCgpZhuaI9hvvAUahVXajeBVCINELyhPUelqH/+NAt+jp3A02DcJjpH5LsZBXbdLPK7ffWQ
GkksgUunDZbiCTCYiRUACGjY51LndFU6Vr12XNv+Ej3Ya8YD5Ks0u+hjabfjeF+3XViF6Yn6ETBE
C/BM9zOvpm7oYbZbiXUxc8R/LM30vd2huuIVDWe/Bsc3KwYvUudbM5NRrqcVvAQymtyFI380l1Y4
ih0lMU64Kp3+5h3EmNez/A2lao2eSHthaqjAK7FAaKIurcdeXM/S0TtXPvnDuq+iS33xSGIUckId
+yvZXzxjfudohWRMpvJLr6fRKBs5SUwztibw1u1xwg1AJanjIFSH3+49pJ7oW0Sv07IpYRWFYxbE
95RxW3ZT5AY0r090DCJEpJWX0Jlf2K21BRAcvvdKp53L2fJ4bArGHK8rt60JwdEsDk4Ggvj4CnT3
CkfUjO7IMcZ1Jptef+vAq28NuZG++9WCGBjwXSeIiS5qAlom3XBKYdcOksDqxjR+9lJtvDh5aZo9
zhmqp880/HQhi2yLbEcsNgBj3crrQBMsVVOE/Ul25IF4Vx3Faep5HXvAIDI3Ff/E/ajoSlF+SPSp
BM0I/PGrE1Eh1oWWf6X/F5ychv71hGvcXIL42DD9JbA/XnvII483gdxvYHMBzlUG1bRatW8RD5sY
FEskiPtQtpsGmmeZTNJJLsyZElL/LNQ5gEj5QeBgZehjvYXtSE56ihA3FqJmrpmx5zkXn3ehaZtw
12o1Aqfbp8WgJv6ARP5eJG6zzR+yVk6kgs9aKNTrZhVcRl8Z8w4iPUfgXs72WUlAGomTs5ys2geJ
Nx1uaMC1fIOA2ZI5I8phCH/RtreKXKw7G8B6nEXIsL8n+5j18Lt23l147+cPyVUxkzWj2G4iCY0V
ZiC+HokmknVK7TFKVBg8ja2AJWw3GRC6/BPcyBjHTNPs5ipV2eK/jS0Gng/klZ2CB1V5gU7+6Wqn
Y1knAbBfrhXmf1btDXXsG1/g/oiq2C46k2Yv3In2/MAP3UROO3Y2BufeLVjQQheHLYHa0FKjdDop
8CkJO66VIifh72WC6yE6mHtEZJTjHyBb9L92v0t7gHYCy+Bi6OGYKCsY/RcPUnv3JUMBsRDsVNrr
DKBByVmL7WwyuSjz2bjKo2xe3jHQmA0/1HtJcJoj35XMtsXFq3msgmNScj5X7CalqsDIfyzCahgf
xSgsG2KfyxLqTJZx6K1DGiWLQ8ArtZDR0zSkjpw+U9ETNmuRWaGTypAirxurUv0KxFb+3GjcNhdp
ujE5ZmPjnWFYiiY106x26gv5hYlc74W5CzfTJwOfwjWjk10TlnSR1tgqMmc/bbOAgYO76e4+c6EL
DQD6EU8+rtGdbSyj4Hr+zBNlqdLzMxrYyoeVtiMfAB7b7nZeIzxzw00cqEwnAX4EBqb3jx3+m9yZ
0RgYyd4Yr0PHXVrIlsGctOs7pTZ2PTxC1/fLTTbtyafs1Lk96sOsyLD6BBp/8n773kPzA3yCTK+g
Le14XREMynOuQgwhNdraTBT75cpvoz0Ymps7Jnyy7Jd7NEAh8l3Cum5ylfXp9ZIpPW1a0VTIlVCA
aniqm7ZSdJWbn553vQfQ8GX7XPNmXEosNgTXv9gWpsRb78tHYTYnFGvuqI/Doc2woxRek1b34P8x
aL6Q67UsfyFG36I4LDiOJLfYM2aUIGhPD/vyeKS+OoW5JdQ4/DeOTN2GY73MKvot61dwJ5Sypr1O
roaWDbUQ18mK8pl46mI2mDp+f1V2GTbyI9Zvgl/l7FZUPlwiTD3ooNI2+ZjKJur9uwTfrZcPD+xQ
pcp1c7gzvVBdMCV8s3nUhx57zNEMsXfbcXHb2xwAKcv5Y2Lg+/jJG2Aq85CQuYzVKg3O2vsnLUcK
C8QUmH1yQaHVw2UFWMnHZipuz1BQ0FQIqyEAlwomBI9gbi+k+nc3GRyYjJPKyuybP+E6//kQ8BvS
hXEuBf8gYkbn8fl7mmO9ozHEdubf/3ODnK7skihVuFNAL0ZdHDgUnMf0CtLBo0wXUBxONrmU5Skk
JK4Cy1hgRhqdexpyyPYt0y1dWsl75V7HYZsRuF+EZBptLtyafzvVVvcWyuZOiu+2vRJLeEdX6OQN
LPG2AhmhL4IQteLA5zsZE1noLfw5uzwDR4afCgHNnO/Jj9bpa1slJfEdvv31JpLGKqqWU39zNYXr
6mQ0EzOC+CDo3HSIaRov03ca+hRvbbh3yji3yaqwoBcq6TsubQ13lW4gk/Gw0rQdPJ1O+UO5l1qs
MGJvkjTWEq0pjUC7GIHmvOCFW83qZ56j4uiKldTFZlEqlIgZvRwPPVhepxmUYjulc9VKBQQ3A06i
NLL5EKhOzi4Lp9Y4rPpt2QEGBwTfgFMIU12plBF0Z88/7UkBLsRobdjpsa0vzVM2Iug2fXHzNgCP
3S/+4zUTvmtnaxnIoKwUF2U/zUm3IF2eePvLu0CwVGZvIWAg4+ucqU07mzzhXOofjtVcK4yLZ/Ri
nzrEsZnyRDPe242TH1fm9AJZx50FlKedWr/U8gHOHifmA4qPCnmr2qMawNHnDwUHh5TbilsG+L5l
G84PNu0XO3tniIAt/ONa8t3seirSBrhh1cocxcnIPY9dyMA9PdDBkvonN4JHo+/TQOBk2dmD/31p
M40lzRncBsafEL3BXVsIBb05TtyUAaSz1Vx8cHMvPkmpbVn1TgnsBGkvgnVqTvbn7Qe6VpLv6aOd
3H1ybIuYe7u4kM0g631rRgtc6fnbaV9qL5Bk4vvQgn4MpxYKLfuPNI5UsWINCV6YfPlluLmqbL11
h4R7Xwul8WebNMMZ8wXKCiJpLWQ6bsU6ztaTPmdbd1vmGiAK0ewmtfgNw9n5TnDI9HZAF2H6k2Ps
sjLpy5pGEGQGvytubJJQ8ZvgD8GBkxywShNrwpPP55+oMkOvG9IQQY3Z0ySHzg85MTAGxTcLFJ46
tZ67wRIOaeIxhQYiLlQ5sU6xKOr2Ca9znYPVGsQDPy8jCjEFdE0EviBKn5nmooMkL9oiKYKcI97r
DXe5YV0PNb3vZPxkceDFMYIBsLE1d7+ya9ii2Mx0KKWU7/8gFXc49vlTPK9UuZm/3GgeaX8Qdq9/
gbU5q4Q7LWIhYsoo9jeitfYZ0KC4UxqiR/YsHvB7oEGsPM4s4TETCg8qYWUM6Ckw2/oUs+SZeBAh
kocH76k+kH8X4H2BeB4yyFjXzluW6hvOAfrNLInAUHlWMPVe6CnyP++W9I6D9KUMYehW4yteR2si
QQVQ76WMUgIsrT7X4akXHg+KUiIX1lnI0IwYbjc4qQmx8Tz9x9Hm2A16e+n58e0THE2sR6VqUtud
wKT0Ev4UUnQxzsjNBDy92CMBI0CHyICF2pDQlasmSy4hRu2NQXqoXA814bcP538dB+NlGkjG+pij
74Sdxu5qoyVJvk33/rvbE1M+aaiLrEBkICR1c7nI6YRdMProu/1ds1EO1KgRCUsH1IRHc8D29Sbz
O6tAsCSZmqkV56SpM6kxBnuxtvIJQCvwjgP0wxsI4//KMXo1ySUyLawLCQ1pQ5aK6kJem+E2rU7K
CPNWYbidYtXbPW2Q7H4PpiIKrcQrNDQ6xRZMVOb3dH5D5lbeDzHRmZLWLR8RGsUEQK+P3B8y+b2I
HSWcb3Z5IXpfazudSsfp8rMQ36ggYsbqgQ+sQLocZIaaJEqnXvVMjbDkshHjZH87NfNpziAYam32
4bO6jU7uKzQWU+EgjR8REYxNMqvMrNhtn7FQDHzq3XXry2/xmufyZwP1Nk/dNgcJnhteOJQtNhbk
5EZgX0e0XL++sszOwMookmWly+9WIrhVavgE2+5qCWZOUVmAsYaE/z+6mqgVuH0nHbyEuxP2t32b
oB9Sa4hIZAjIKSYAfr/5R/TZETKNCPlp3b4sFIMqxy4KCK6ey57fjRel3hElMjNe9tEpopyYjXH4
4ZAraNf1CWcUb48+KAaM/oRNEAgzwWsAhODzTs+zG/lCVYBMLRCoVJXCJOLXHqWKKp0Gi2BirkYN
kLZpqFuWL9hCcSquX2UlKxSQNjP+S0Vq9HVjbFFJMak39oFMoQAlc7jZXjcjmlc6UIZ1gTyQgPYb
aAtRHvWznB0HbP5wwuSLxBCjg3zAxPGuWfp1LRLMKS+PFcRKTY4N57REmkae3acN2Vq/udRruzJU
kOvTZkLQnyNIVLLy7tBJR/6B7slYv1uG8GSXucfJrZhymurfpjjYXlKUK58Rdsz2KD+85AE6+Jdp
3qEJZzde5A5OqkCVScekcHjFGdg5/izGifHggjMPIUAx7mtEijnjaDSfX8i1Knf2LBzKdtSNnVZt
N/5c/Ml+Rpt2lN/bryqFgGqOYk27cDBni484f/7iKN0W+vbrjbCF4dKjVzbFxAQAb60w8gTVfvny
AdOi/jK/SayIEARCMakdu7hLoHTHAFE3Uw4etLJG5w4s58abl+N5nVmRX406ZxfWb/keERq7Tq/T
wPemAPEVD0cFAZziLXFBRhaa4l3rGY6aUwiL6FNoO8Nlf34KKhX9gIqMUbrg8TyaWcXzntBI0mhF
idGFXjehnle5V40tYwzKAxnU8DiM/398QUS/zCMF9pV43ueqngc5iXMOOxHiCwDAnKQ2fy1/AiVg
U9Q3XSKz4G1pTfVpSogmmw3qHdANN9CYRrgOqxUQfdzqP7NlDlHEJ44+wCXtQ5u7llV7gR1fHwcB
m5ctm/H2iWtPUKB+A6EJP8B4a8PQGZl7hCRHTygf/OPFM/ns/EuF8EPrccCQvGUbyIHY7v1kj7a4
fGBd4KI9ynmc0zrTkbmHDcw1AaW6yHNM/X3HaBZdqKGuE3nw5MahM02gc+jzM9O1zl2WiasdG7am
9pqKemFxh1hz3SPvpphWeQ+jZ6d3T9vzUHTXUfB1dzuUXkejxUYiQ+LHAqumWx/lDaPNCZNOzr86
QadZA3VkOdMsPUafuxSZzoYZM4Tl8EKwLjz7mW+8juE0a3pjMTv87kFAYeNxa4wAmAX1eS0T1MoG
diXDmktG3UCPgPC3HxgywuFjQMJqp7dSJE7GYc2deKsXP0Y1lwZcmgk5S1y5M1KTg3OowLAUCOjB
r79djwuPkFfgeZs+bcZw0wmBJgyhAccIiK27jjOMikg0eNh9xyb+3vwTfxpAN6rm45UoxNhWZFfQ
J1qp8pltx85pFusQl68BFd5QDi0nAaNP8Y7mSlooqLt6GMiGYUZEwrYTSMA6fZfsXF9blaA3RLGo
g7+RgoESl6w1nLOHdejiyCwdWdkiqEwWs0mssWo8wk5zOb43K8Op2ZuL1+8YD6b8cC0zkc/Ra9Ng
KiGqQ150qD+lJxSZmepttyEJlL3Y+butt6SEg1HI+trG41aCn5OyqKCStQfUZt6ewXCgzYbD+AXq
6XwWy2+AMtUcY7Tpn1m9DQ6IZl/ljVPSL+lOoiwDYFz8WfLc+AXZGxPjqOFDTCn2Ht5THa4wUu65
a+8jkIgx4FkHtELBmR2KUkRp4Li/2CsQbvjC4HD/axQUfzbBnIivAJCWor7oaXV7oub3W/tbt7Ov
7WwmydACAupsbqyxzPoYJB7jqT+8ZWiiGfpfWi83fMl2UFFMb4mpf565zQCFsfq7nhXXzlDrSU4N
y1qLsN1h+Rfox7QDqkiivLvxVeZPyyZPQ9mv92mudyDK/6bruMehTA6kpPFuf9kvh7IpzQ1RxLa5
YEkHSJJVgL/e3FMzqCEvpgsCt0am7Z09Wk3iYSDkMkCl4aC7RK/zogNpYFk/faBlAnv9cyszfZ8g
V+SvLrLyVnF+hdjr9AZ7xEvO3eAZzERsh+Zu/9PaHSomndFIVuNS3mu5A+zIWudUOzJk33Sc30d1
KiEsK2n6ebTeFPxUeHl3GM/eHpUFi4sy4hEsr+hFXwGS6n2YF6PnrmQjG4BnTUIJ9PKk84Jw8R1A
pV/UatHfaFRQejvGlnCA3lFXNNFxzqw7N73xkuyUoA0DJMDwPnQwfwjeAc3Die4ycDYIkjmClLEA
bpVHRpg2lQVSYY9uy5hgZHTOneRhJiyVZacUpm1m8D/GaT44jVnXOhe4yn+56zYX460CIGlAqu5m
aoQfvPOkPo29xhjbzB8fXtnGb1V+OdKb5/wffCiuLcqFRJBqGaA4fqeKuPxA2Sf3Fzj7pxRdnpEk
Sn7J6tbU1lwyVT7M2+X0j4PX60ySthsC8XqTY0pIzPSSz1Iec4saWXtd6+aBN+Y4d7YWdk8fflcl
jQn0YVUXofjMeQfM9g5VTx1W20+I8Ve59i3VN7jFcQJtlDaO94aVU7xdvvt/8utXHHQWpTzphexS
lU6MHnZDh/LcensZdvPs4jexE0vZWiTMmGYS2s8O99StVzXEp3tS6aLY6TWt0ARvmKO/QA+oZZfP
hTHXvYR4aEWxbkFxgiMwLNxrh5nd9P5R1jhSUDQA3sqc/2tnYSSZYZ0Djt7ordCPSZDlWy1Ye0qB
WjrCxl3qLCQj73zonodC/QKVYp1bPMM3o4gvBMflwa+omfg6Ydp1QulvKChYGjrbMSb3sXRVt9Lh
GLNCR4G6UWTgaaFZqZWrbTnsCp2nGkVdhUsB9/lrkmpbd1UcpIUYddzCPETuXvCpOWOGV/PUuytj
Qg+BSXdjSyCDFMsCsb6rAF8vb05yzfOyySAwZNPxkmhbkHB0buLMC55m4AmE5s/WYV6Cw/9fNod5
ga2FbOQz1YGxt4MkCH+VurL7Pemmj0djR/id+r/uCjj4kkWOAcwFAC2wqXVIhdWYSH4C5aDmZGKx
GUofvv8IuAFms4k6w8JJQyttJ1dL9KOTSOtLn+ORLmWVDmiohf2sfFW74t0N7p+kad+7jPNZIMb/
f4F7fQqxtE5UWoPCoLnOAC+l65/BVqGd8w7lLvZ4OAx29I3ipBSmlIhDp/a2ylnYZKqiU3Q8y4GC
lr7B6NlL1DLc/s1L5c2+TSFhK8UTzc+AD+GARnvnNx60RMhFyriQpa7gxo0mF+BZ7aiRHMDGYZTc
QTn3YOmE34R8rPKbue77QXt9zaacbueaZzyUPtWfINYt4Uo+zv3UoAYlWAYFNcm/lMHpLRHUrlf0
EY2nnEEwH9xz8e6n9IaGbplCwo7x4Y5vzk9doepq1mNSIZMEg1WBk0634Zh9nlReBMsgNu2UStSD
hDSsV97hmwF3Z71Isax+VyJcTI5wDT0djiUCRziE3n2UhjxNiqBW5teTAHWTg98ch2sQOoELzdJQ
7w9hYtxofR5Ex8j2VggdWpYr4wO47w7jhAczQfvMQgL9TCwXgI6GHl3MKz7zuhfO2SyFSmH/KhL4
RFgobpCK2g4ave61nAEsc1PbvVKFsR6wofJK4U543IPAhuXpQg0uFgNajNDwX/wHs/s9mgFfVCdu
s0kfA2wayxxvpZGuHGUkc7/PQA5ePCaRB0A6cPqP8cjQ41VvKCZGSjEfWtuDE6M96kbksazWuVV7
5vxwQXEuwTfXllI0GfAUou7AlgDCb/FI2/6oBDoyFYl2LX3v1aUESu8B+7iwB03aiSDJopxyTgDJ
R0aDJF395Q8pQFCMhSHGzemd0mZhoujApEaA8V6bzkJV7ZtLzoZQyow8Zj4Av2dlMeFF+e36YJ6l
s/rLY2n60iqZRnWfRQ5m6+ch052vXAVloHHaK6ZrhQ3Ue0jFtBjAbcGP/bXsE6B9rRWGTqLabJve
ckn3W+kXvoztKX9xfVEivY+h7sVqqMM0lV+uIWWs/j7WAW2isN1aZEwPzxfTem7a2zeArQ5XrFBK
kIPslb4cRQ2Yar2NIaiXxaWp20ewEQLSS8tmLJugX32QPdgqM/ExoEJFk16jY3pQIMNbPDYTNjbN
IFjjkxoWbK7TABNHy5xiKEJtc8IRIb5EvkRMmJQ1QysylGds1q81MPI6UcBai9bC0yWfG7wj/VNq
skXCqsO+IX2FVXVp8+2deaxSGbQIWHdn8evw1iaGnhdkaPcTnqgqkJUbjE6SW7YXmP+n0niylY1d
DcAO7AztYhEj4F861q47w7NY2ZIXP5VORe5Tag3zrsrtpEqIpArEy1DxxDEVr7Dkzt8b+iu94qZx
lHcrVKw4o2iwOOEdMOlktiRBX7P7OtoHNGO3pEEdEq5+Q5bQnwUY0Sofyw7al89GEHRpRrVsLKIs
4LGzzQz6xU0uz73xEF4nfjTSghBzwxVBpjedv37Sj3PaKUgwbGjYllMAidAKA8bCvix7eNSoPrHR
UaOqmLQxbBYfBJXsVfSGSZPeq5S4Sl1FBvRjxWtkH0xUW8/IxLKrXEr2QUjy0Dj20k1moioVKBzi
uAcKLOPWw9huFVqUlqwEOdgl7/Bko2Yoism8Osne7Ea0pBmxzbmPzCfe9e62DdUCPM/n+dF2pJmb
OMceOfoP9mF03gZC1pBb6E9jYSFIKjtZDkMLCgUki/TekHwnN3HrpLaSCQ5y3+oJpcGExSoK1EiB
HVFAB1n1VGvTCVhUIifIhLB7/8UHQ68EH5oVuWytilCtF+NVLzijMZiQ37J/P22pvmv3+LW19twE
5zINONp257X9v3HDdKe51iREZpRDdXw0LNeKRvsCC4PzVWvf/Zow896TUSWv7XO70svmymQ8Nvqi
fFj+F3B2j0vHm1wcdzlp7Iq6BX3AnnpT1QlifyVXcUibju3fvTCefOm99f1hzwnTFNaAG44gLbeo
n1zWkYMPY89fbLTZFSeasgpqHjhxdfXKbJd2mED6Xd6igarzBv9Cz+5cS9qZ66XHSahxDdpQfezv
VHeeQ2m/uQgBJAPHVgW6f74Et+8rWMf3qj9rF8VamyWWK48AD9b2TCcvrUs4MDOG3HuO7eopcUqb
KC8H1cY9LQREHL1ZqJtRhID5q6Vu4mKr3Pmid5+v74choUK52yGpotGJYhcJ80BN+ZQAuzks27rO
w4CUrYAFwG8ukmX0VuE03w+qwwWY8/eUjCGBQikQglmbbzwlk56XTpgIYKLAnJe/nJ4+OcqRuRLx
q9OMnZ8fNmgfyOOEuIvk1UZRSL2F92ERX4u+HKg8BmuwwsXbapM4UViJvUcOomcQKAyMiW65TfrQ
komlExSO862fRLTt1Cp3+KOrDOJgN/1Z+izKRmkG6/9FP7SkUUBh9+ZolSVtjBxLwmjfagpeUUns
+oF7tOim9gnJ19VlYqLz+XnNqGB1rq9RyvH+RIJsVroGWO/x8xH1kr2iCyhKGsTKWpC3nqNBinUl
f17KTsm6uo7niwYpBQAH6iU0e8ty3otKWL8CxOa2CkE9Jtg7OQMNZc8SuKCd3Zj9NPskvC2CXAM0
ziLTHq8x8X8Jy3ECBIgIwPstGsKy+Ztd7H5W6mFxm30c4aAVbSydCQwbKMhcz8gB6rSPAxSzidsH
MW2M/93+SMFRYy6+WA4nh+mjguQbSNcfyAL3TeGqZIPeKK8fQblFbMjmKqXK0NOSQli3atBqokoB
bpZyMunMei2PFhO3lzsxqi/tOFd01zmJ8vYMpAqhmrn49lUlAhorzRW4Z0Olnb1uUmF7XsS+Ywuj
9uFHVPEKnZUzB/LEzY28oturcGjHZRjyDVzu95yMIfoc87qnXvDmAGs0uA6nnfKVM7XYW4kcCbQi
C5v8SGK6Mah+mVf5feDoWZEKqaY+gKhpDvpSwgqRcpTiFMTyUkoqn4oMfo4ZnoBtwXysCJNpgVTT
LiFNCLVTsduUjUqh9mbxeHWyLIxd24396IvUEcE2fTr9/XbUh7VjTrnWiiXw/tK8zr8v//ACCxlO
VYkQlJaXNNM9Fr8OEh7Rv2yTcj3s/XXyXlpvGWnv48ofP9NK5BntvTu4mfpWKeINVGNZ07g8FcAl
yGk22oj8yQz/lw576stKaIyf7ba5+0p4dIfeRL/5o02HeJEUj+LdiPc/FjldmB/9IajlN3tHARYf
p0IPI7ACnsq01pAt9FsWVOWtf/wy0iUTgeH065VSrhjWdZ6nWTxyCsB80nGyiV5YfdQIDrDdfM49
d83SNl/4DR+CnxvqrWIlmw+r3gYUwW5WdPoFJOV7MS6ZYHgVvfrW9vGPfm8C0L4TptBurZjxmqVJ
XDLKlSTGAtE2GGsMEIjuctrEzrPrPRbPjsSELMcEXqr7aR0NjTmuYKfymGxFKUM7O49rGsWoRK/c
tJJ7+aQv1IUk2Du7rSLDdKgjjzq4gPutRwTpk0dEvgTJeS0HkyujqxpGIfpddatE8edL5oPURbs6
ydyAq7pDjHCoBFJM3dxllcALxrVRv8RigE1Uh8kCxqcPP1RwhIunE0li/bm87Y8rfHGY2EG25nRk
qPYvMgS3GFN4gLpIYBElT8EbfwzjryjGr32J/JMRV8AMvujjN//bBZNvJkBMRgXnnZur8pXAEZ5w
fuK1SA6ZYYDDLU+SX2E4QbSc36/qrRFAM2rvAjfZyLsNs1a/qGcZwFcmAHVEW2ZCvEfd+gyhIv0w
+NImKQaaafXMVYBgyU47tZyKlt3HJYmAHNxaqoSfSYoLnxqgAmquEP2C2w+EthrXdg1VbWaz8mXL
1D8K9ek75ykJ/LZSKRU6ToSHYlMOXUOqowuOpYd0kjAtmeFJr3PyIuuOeWtaqbhbhjIyyqmYDncY
ZxNtglRFqpYVpDG1d+1f6E0jer3nZGypK4fsDLJQW29qA3TvkMvgf+EGPWGhmgOZROxwymIhhHgX
QQBjhqB2FAVn7gnNeEKxS5dEWSn0T1fp/sdKWWTXGrxdFL1Vc4ukGepdkYG+p7lm2sGhH89JaxBz
dcOpD0mkIbB58qr/qnPdc8+XS0dAFLWQUbt0OJNZ1WAp5A7WcRqAwIVr0m6fWxb9Sw66uwzkgyH0
MEd0ErmzBINpG1pvNiQ3qsEAi453p7htBqbrRBxi8zWUnkADoc6WiJ+lqhpQdLy+8HU+w6CHUvCL
062B4E2ZA4zY2CB7tJG9XFGPrA0yzCK5ZMRxMGNaH8giHsnPVED+ouRW3jtfciy39YImbf2IsUJU
j/Y80048vXcXB7VuASEa56sabTbPSHm25GW4hQ3hEAvXhPTv1gLty7APL8fsdxMvlyC7MogFUr1i
LewloKe1rKGuIrZ/W5CXSR5xU7lCv79Ok9Fabjy3tOTJo+lVjertYuViMWvvTCyWuWK1tj9OWVlJ
ZfReY69p8Rsj1zZ/IcFOCOc/ZlE3vQXaZIas26oAh0+QNXTzI/HpW4Wu48F+olADnb6rpuAcqBaP
34TpsnpIAcumZEb+3jy1W+r/yFg1OzWb5C47DyDrfuMobAtysAuPo/i04HfT83alTeTq5KTz7zX5
g4QvHkZb0FRbjxICXS5mgZJ0w+5wEqf5aKJLZyoWCsU/KDyA/Zma/T1Po+n90tgWs/C5Pu9L6PwJ
ZK+a2WMx3/PmXmxGtv4k7S6PdsyBbQcDogG9IWufVkeUQ9379S+fmlNw4q5Uy137+VAxVXJdNBVf
x8IRnwYLh+gTpgczT9owELzVwMel7XbF9ZNaRhDNhgU05hLOARnN/ZgvqxL/m7VhNtUJCQd9DLD9
iLUm8QxSlimAbzPWVx7Qp+7Uab4n3s4OHEeQmjhBWsdwEtOw8ALwDROSgltUhWFNaQ7A2aSm45Hw
qbZS7OVcNJqPrkZgjxJVT8IovT1tRK7JDrPnvZyjAFyrObCZXvkSeMp7gtJKhh2UxST41kTKwVZO
5NOeyFqcfj9N+WXZpBAMi2EMUm5pV5V8xqTU07w/wXi4ZLseV/cvUxXEfwJKzebEZ/hQX+3vUvRF
BqZHrBgnU3g4vKwK8lKYgS54q0v5V+fsl43F6RfEOshY/J1hP/warn+nImM1EF+QOMrBCstGGCU1
F6TOypyLW9/hOLaQfdQ8QeAAvlnkPcWG/o37doVaomKiYap9sSJUUXDyq1UfbekEe7GiRVl3MLN0
9wW5YaKC9V15I10sCptnvTpWkArFggwzEt9J/HfYv6oRessYiCiv9RsGtOTdGyjQZTG6yTCWfgyX
/md5bMO19ixumk0dFPOJ4/fqdzbDbSjXJM3TGDp1dOwdviEOmH4MDFakrkxgMEAtx3/qDLaOB1Nu
z91Qjj+9x+hsyFtxg3rRsELkNORxmaugLh2al+u92EuPim9VfROai0AeyNmKY/hvDa8ENI46sRlK
Ch+a+Wp5bcogsFA4oScyFjKofKrI22SuUi9iTY+8AFmu9hCDK7/kgdmvDZmArGPAcWRxn+m387N8
KJ6FsErAO8JnOeteKD97XgKLW0Q8ZQrjR9geEG+PZZCLNPkux2ezRp1V7Tz4+fCU28pT9rQ4GShK
wRYnUiL9OtLm9fW8eZJWYzJdXZqf+rCCBM1i8kgW8gjOFU7ojVYqmd4pRBBiBk9qPVTzfmVt/Yp4
e6/PFmcU4kHQ1aXgjvA6ALqJGvGHIYieBBYHTVHrxTmcZpYEcw/IdJLhTb6cAMJEnZs6yqdykaPg
APltB8cKFTmWn+YeSPjcmxIoPIAKdDKxfXKkBDirjE+dcGK/kXfRkeYrwS6ULGIiRY43HvchoqyA
FDyCyxA6SvvVnXG9wYz8GE9VeIzHM+VOs0mjr7bBXCJq3cf9Pectp1pg21jDJgLCv7u8cxqr2i/w
awAJHwYQwwF8MRAiLSvEHH/dXara7jzPwTZKOfiM3U2oMcfXTKwRLOsTHNgukSn4BLwlv74FkTWz
nlqvFyFrKzgTkCLvoHkWWfUmFsoGtE4FO8f3ktE5YxWqOBX6Rq0HKt8ocQdwJeFMtX5dReJ3F2nb
EI/VnC8vz2bm+De17AL0MKpEu4sjghsQbWS/1PXzACLWeXufsq1hXrYfz2P4uWPpkUevhGEGsnta
A3cz/QjmZoxFw4bg0w6WU/e3VZb9PasjwNDMGdIuNWQcAwsgFyK/XjBm2ZcxNgJ+I2oDFHaDgzvP
e2F++iZpYaY2yCdW2sDXxNRhAURJ5//2Mp6eEKGf2SuYv4j9CYvx9Cw2OKAk19MjWQP38JSTeftF
3sOifd44tCw9ufTiL6j+DYDuFg5AWuFdAIbr9Npbc8ylqFXcHVa/J+Bsv4JT8JlE8uFGLyicE2bi
x+DotuSCGmcImi2tJoD0byj6nn9VEjTczuy6XMUvimSIfV5qrYBiMQNHObgKq6IM+PXtbWF04ZQn
cqsDq+u2jGcnT57sBXXxlbzyHtahI+BbdTRfohEZxEYBKIK52kJ8myoWXxScvRRJNydVhzY7Xy1d
wMeczalcnQ9TCFgr0Rvl/cUhoV8aVYuZTFbICsoDzalwP6i/HowXCBIv6fL6ZcZh9AzdmfMXeJxf
hVjSLjOCFdZQGKQHK1Ely40Nmm4cx4jsOngZIjQmRRGjTiUVgHYOrMN4N3aqcKFJLj3HDUZkwOTL
v9bvH2gZf/1nmA3TqgCxOM8R5p4bThK/MAWsjOzDR/CqXZFphsuW+s3t6XqiRR1TyShj+vu4Usg3
7o1nFt/QPVp5UlPdaqOQQ4hHsG9F4cDH786W1sQA0Smjm7ZJm7zxiRY9MTZWtvcDv0q3myUmnaa7
jIzWzQIqTnw5eXcxOmCDGEJprMAD3KzEVmObGjCgRYXVVzq7GuJv5PNpt611vTuHTpBjvnydROyE
DeHSoIkAWqYM58DvDctPqe2702jM0jdBh/dAblbkZLEwqK+Tz7gXmUs3DohdXLanpbgOgRGg97uy
qmRQ2s1Wb3fVphhhA2ecSPYXsBBO+j1dIgs0+B5IHpjVx9h37OPYJh3GA2fPVpXykkB2nordGthE
uxZPp5ocSwgTsTXLOxXl8QpL++g5QTG5cnROIjSSgmnq2Z4eFtG0Ij4ql9FppoW77juEWRdy3SMx
hVY1IfLeA73YE1yf/G7nbe/tjbbXOVk9SMZReApfGpOXDlYCxfsYzqZsJZhL7GRJcwdn3Hgp/f3I
X/+BIHKgVzmwahqmHDmOKYz0ufYBYRDhVQaSLDfOVI7X4tflDLbZWrZCCgWiNPKEx1lGAMUndJKV
/hshrl9L3FnP5Rpb5jMZ1r3YvvQUMrdCQMFp3+XV4/VwygYukcKeIQAwudErAKCgS4P7fbE+MS1L
RlXmRfFR+UVym9EQd6vH4lD9I9ALd2DDU4m3rHCdGkLQbRmqsdudFBoMeVg8zpUNmwh9mQcDSO1H
Mx9RIhE/CZ/SeFJu3fkjRwhzcx5OS4xVp9/Rq/x+X+kv9GXdXasJMQrLRpFs4wHzDEhtVa686Q8M
uYx+Kxp+GLfRYS9gkzaUkJLZg1e72jal5aJ6tQ8Ac5bkReMPTrc055ZiObCXxrzCnNinfvN6jt5l
Y1FaONq2M7cDy5HIfE9AkJ+nl4vbI0bF1btVroS3x4ACqr2EjZ0ZV4n3XXtKU14Q75viDREY5g7F
CJwth82rKiCT5lKmxPdWS6uRwGMWP7YV4yfiOpmIzNucyhSeNW3qKqOvFyHnay9EfmhqKIt+bd0+
3PXNyMR4TUu4zq+RjDrowVx6uj9QTZJT/1FAs2SIUncJbBZvU0J9FnseA2/bYfrE+kR6qpnoCg84
6SV3DW4PQk6P3pLFUvhCkO7LWSOxG9/av+Q3aR++4qQGpXwiVYMWB3gFGt0VjJYXaAkE4EJGWb6g
1ZEJXiq6n9AljtM+fgqjRBEPzZZsMyDdbTnumHXmuaVtc0t8NsbZ3Q3BzII78Y/sL8BOJ8me7VD5
z1aQQxs8EmM5aViyY02OMWw0gnqZash/SKR9WdOneyV5aJvO3jfhaj3EjljzVJEm0BYRYFUDXl7j
2R2f+VWli09TOJnwRIqzoIDWnedYqrTG1X/+b2vRn33KuSik8a7eb4MfAp5GISC3DX19yfQuixGY
vGNoVz6jEpZpR9NgA9+ONwF2cR9nf6uzBWYNNtYipvCyk/Cu+0asm4rNPiIgg3/ng3xRPUi6eFRE
6asqD6OIoBL7OJzjNdEJHhf3s81WpZa9WlBnHrxvO1i/AVr2ZzQTrl7f4D76pHbbzbDfXW7D5b1M
Sm329S/VCzV7wEdRefyCtwC1637Ssi+c0tStvgRBn1DfdIQlxZeXH1tUQvy6d/NEYMDryBnAnR0C
dvGZJkKGp/kh7IfLA0LlgHLXAePlchbtqgGUVLyG9jcfzfeZ5qZboa43mtjuf7ol+fAPmEPCVjDI
ANrU1YkzxhAjWYUQn96Bplf7umfbJURMHPbvbq+oXeeoDSl6cOotjcLt+5O32M7mrHV9WamMIhwU
6Dzc5+kRRrUcyZ5KjccUvpd+hmzjhKJGb9C8GVl3hdUk/v+ehL3qXBYBOseMSEhKRWFjVaf1qqBG
KY93w+y/iUaRnGxJdWtMxTBcVPZvHAeD0XTireYHb4V9vOgmZpsjjlWUNvzXFOX+Wscr2WBEN3zp
XJhO+mhsJ1PanL5IJDEHpdlqKtICpJbSBHF7Apxzmf0rGoGhkQlbfwi0sPZOSBNbLWujVdFgpECj
G8A7XDEVP4LlxVIJsZMY81lGXtlEE77p2KH/o76g31+sy2xWr1T9wHvGZaHDsU9LdiPlk0YbZIbL
nCMDCJyxhDkKNC6RBZTYlF9N5RBSn1DPxxAH/7LGCDwqd7aiSe2fz2XkHS2khIm8H2+r4JgU/f1W
tnnu8jo2hpZsOvigIn4l5pS06sp69M/BtOiLvG2x2/LRZr8rXi3xsrxNhtZECBjh27z49a5g4HyX
qL+yzOmFd70yjBKkhAyW9eDFZuc9GNtLRDp1a9HtptRlDYaC472H4Rdq4iREV7HePUiVaq4bxIiT
Rw00iJUDrOxPWbPHfH+glN2lAz8ijnlzhH0x6baDZ1XZFDkHp3p6Gco8kUkU2eultNTR3fob73GT
l1cPvRZx0TrC3ClnFjIzx1MUrJKNg4W2FkYI7b/I/5xZim6WIO9TQ8TSDpCwQcsUHL5ZXViX4NfA
HKO9/E2XvqQv/wz1h3aod9RThcf4qBOIh2AzNbRSo2J1jAGAHbhrSrY0G0QR5WpB0THIO4ZW2E1O
IhOZS4/j6mrvsUQ4gcE5g0sa7HMCiVKLTgrEQvtXiWokVcJH8aHr1eD0mHx5WcvyJPL8E61twQog
rH1ZArbd4SBKuAm/oMoJHRP3W8nhK1BdwpHdV8F1IrDdi7LP6Yh/woPSOeuFHpJa3sS2qkzgCrUU
jPn4MsdsJgRskCY6LZ3sCBeobSGshasAFkdQ51PyTAXv4U/sonmzR6+IXRnNkAtQilsf3DmgSFbx
+obnFw/Yk7SWGMEK7w88FHI5b/5e9OLzaxOyEZxOjOLhaJldnWhfkp24BT8mW9Nxa2S6ih1gnPko
eVln5a5Zz7ZqNLU97bkD8TCm8IZ04SKc2EJ4Ak3fqetHx4aNQgQO1dxlQa/JP4w9JcslFETdtB+0
o6gdl9AGdd9Hhvh9Ug6wgGMQN3bYE0R9Ne5o2Rs3mKoq2vUh8cWjlQAd9N1GJlQkFiRn88hM2EJR
x2FsmpPyVpFSIMv4EoSudFClUYbRkXJNfKPPacpbqDBP2TJG9cY9BjjBx+jfLjMeD4WwGLSkOkX4
N5stR7TDaZEXgTQwJmyZ8vxWhCVURMu+QzmutQVrIIo0CF3zU4odhrlGS4N7Gb7gKuyNCvsddUxY
EeYGPzg0VliC7+ujmrd4eqbiI13zbBn6L4ODBbPNPNTRayxOimQcpbfqXM01UlAQ6Pw+DxxTGXY6
3yLc9GN83P0fw6W1f8tprNTHm1xcR4GG9+VqdCiQWSG6ly40ywi4Ndu/pCSVATodPyYl323VKITQ
lqU86Tf3KVk/62eJhIDWF6LJrlontthUVa99LMVNspsWaZzy2r0Q3pwAGs83YAume8DyyA9tuMHx
EPtiIcFqVVHUHwNcQOewzxXvhnbb45/Dp9D3d1HYcTsv+dvmpWHqjhwg6kZk0DLODQiTXgzTNI1g
mgt+Z9F51t0LnDB5Cuh7QDCC2dD3UTuq38xgY1EqNHmy186JMDAniYa5CZd0TIjYaygoqSN2XGi0
195C7Mfp+gCcxmUQ+Ufx9IafTmVjKo9U7cHBGC1zn8OYGxE/PGEplhh9smIN8tYGV0Pmrj8jJ7r0
Q58DMDY3gsXQYzRpDCLftUjR5NDzzSAPvhJB1uUh2mZfDefd1wJsMa5rCUIyIozsz5x80NhURMJr
UlW02S1JaPDWlsnTnQq1Xveqrt2VnjD6vBgeFrH5TB+5AVv9SDZj/flaWeWSmw1JTj95NMceQO2V
+lItfOlFduUrGM9VzTbylXp9JH8G4ziwlam69DhHA93Hv+Hmq8BrjMezIHMvA5x5xbnbHEmJrLTZ
3Rt8sIQFKnk5CvE6y5sX1jnReztBGRYidHkonmyQjfH/X3/djYlTGkwWVt+ph/3VDJ+HoO8swB3j
wbjW2zzlk3bskEd4Bl7AbYiKr3im/keaPYRwYtw7RT4Ei6W6F2WlIJBkzrx2WYftRbSBE9n+MwiT
6DhkQ+tAnqq1gKRdDKoafxzat0Js+fjIPQg4qDqrpV6c9vkQa8EKXo1HCJ/vRtCyCF1KmZLiOJrU
Rl03vNmJw8NunDg8fM68FZTiA4KzZEBUiYTdBKM5T3TL+gWTWjkB5SLeuLkR9Ujgwe4XLk84PPWL
gbQqnXFzSyzOds+/cZsUTr6YT9VJ7pJ+9x/OhP5R1yLs0BFTHzCMhT0L05vzV/+eQEndlO8SW3U7
QC73KHsQrtiLf1Be9U8/PCBbSXpD4zkvgrMDTAqoiHCKnsf8DKSiBNmaDA3XZDH9fV0h4F5k9aS5
IlIIRHeDKhkYTbdl/FGjVC8Gu8+Wqi4fi3v45zfbjHKq+2HIqaQqVln9W5KvX5zxQ4qRFftRHgrv
P+b0Gh81PiPZa8ZfMg/weaJetfdlFUBPoFUcwLPV0LhYProRKM0JNzvSonDfPtE8esGlBJV0uq9j
KzVzaAQ/4XeiJiieOAtBMRsHVTQujxtebAUP9YFZqhSgclN1GIkbs+vM0wRmS9R44NjAlPTuQdof
9Zgi+Ealv+Zzp+uJY7wayqolzfcRYOKrVtscEwPLInqP9wFSb6ESkan4UVP8McmBNMz1bVR8vQ+F
nGubjsx89MV6GZnz1zewWKRiuA7U7XEdHWhI1LBncKyA3n/B6CrKPEMzLVUOHqEkXeNYf9/caPve
Lx2ErgxuX7yTVB8hZmTn0KHdNIFrRKqRsOgRtLLqbTbdXTj3rP2GnW0z6YHrf5TK+njj9hUJ5qHL
wBtDTUC/JkRa1ZKwOkM1zy9SE6d0aTUP7By0CcBMZaFsJIeSgpva804IhsXkCMxf8A6GI2s7tggC
4sxFKXVWjBlMJGQFq7vDd7DjjWxfgKsMAEdQ/bdy/r+ivnhRsZrKOhEuFrV3AayuxXK4CDm6kBCR
O3KkWijNryTe2DVVr8HvuQRvXwdZWACnOTWG/mjJaVy3IcKSTYDEJQio1DbqwSFnRqES8KPa89/Y
K/O74oJWbjR0B/Uyogix32rN8w9RRkHK/ffUwgGQf9fCu2k1qL4p8J5QymTNyg+DrfGntq6l3Avf
AE9TH+pYN1RtP0SQ8IazZVpwGJGoFvS5aH0WQXb8e0V3EuvRIiQpuTWjFPIMbrqLgWS/MJe9Ondm
8cC3cry87yCK7WzfH9Hg9LPlQ/onCfVNMjpJqY+NWCHqSyNQFPF1C3DxPjdDCIf7VNR3y/C8Lnkg
XUAUlwf0vZ7h5kF0gy9hgihpW1c61iksFNDy1qW329O6GmLrCFXxQMSsWBHE99DUT3RAsaWQLlJC
s8e++/GE0veEF56Jb5sQGN60kxrRYj8ZLjNgwrsKbKHOmfAKzXfwpdhK1EgLF7nsK1tKcm+t0N6r
YnKD+PgodwQqwyym86HWi8IXIa+lZzSn4iRCzis1ELZJLRrHWejTM6G0OhbzvwxYayHg1T6dyxDm
o117NlIiRv70E3gAFVdwm7XlTpQqLppTLTi4Es/GsypPu7amD3iJqZcWq9ZdY9Ca6C01ZWef7CGI
rCEE9BlKIRaIS1GTTCuMzs7zSznhKdrn6wTWDl1t+5uhmxsfVlHO0JyektB384ZvSnl9FnW2tEaH
YtoOcdWyWgxQfTEfnOSFEaBUlWp7Md9lRE3nS3js2L8EGcRGIm6burTmm75wqjkJruo8zWNVum8T
1z8FCTUFHtup0f8U/nsQDbPVNEA4D6/aCL8Xn4iLb8Gm363tXuE+Mq+rP2Po7ra3FzvzLFX1E8L1
KwWmqvJ9kQV2ss2ZACL6JFSoXi9WJEZofOUIpkLRrEWRKUO3M00hz1VdiXJPA4zZAaBMK2PBWgzW
2oupEGpNBj+i8H5Ejtf72Ro+rO1oV08uDtjw0y75wtgveNySoMFrtQQvIwSZn7rWrREOrqtF5PES
Hfzu+2PMvSBKAPO/GpOLcLHIfd4v5LTxYHIAjPlCzuyvu+p8I6MXMzLP/Md0BVNhmkPc1Zf/OseG
7oFSVaWiVzq3I3WFXe8qnj0LQ+8/RK54bmEiywUMUIpsxKIYvKNmxpthEtghPdsFx3X0oZx6ZJJQ
GJ2zq+SANMf8MEucPc35q+UiUJa9mXhleM3EUhxESUIpr+p6ULmXLcM1cT0PtPZFi9/1VxUO8bUS
TVdhMn9hP04XcsRuaqZfrl0yfGuYV3rjVeUIEGjswA+58bms+aSiZeCxRQUsSiaFpp1EuRrHPLmB
1S5r/K3QdRKBvtBecb0f8Qh16xAu6eqJNkssIR+ZRTmspJry3XSOb0+qikeS1dK538JaB6t9RtS9
jrwOkaCc0LFhxJkJaMbPh97y5nMyF2734hgOeqWVRD9HKdLP5PZNoSedDs67rCqu1JSqy+lmqCTJ
HUJcVpAgmzG/pjWVtvpgyzfyg7Q43wJlY7uNRUjwOjEvyW04WRfMVBEKIkOlQ2rtJ151IfiGzSvO
ruEmrNlyMwUvMMx+4UpaKPrHjtz2nBbmo/3bfPc4sOpO2XhRQf36VIX163def0PqZ9qz5AZB1gpr
W5Rvp3jP2xnAnP7SltTLdYZW+jq4M02Y8IldhmPdWX8RD8J9fhOUqfO/hJz9a1vGIlkSCO3zpODd
jmW0EZOt+V9YMueOBayGl8fHb+ySXcIVr+MyxNITa4WhM7EWH6/t4EONTKO74MdvSswC66QQxtWs
7i3lVSfyGXInzXiE6vNixfNy22CCshK1a1zSh8IRcJ+nu/J9oqdjNBHkXlvkW58cHJqw7TJe1eQr
EfotY5tvu1Waor0Gn7uIO2aej0RBGexSVMDf8/YHGGzipBLIihZrlvldEOUkrj00k65yjVXk9sSC
LCZEEcfZ0cL/Jadl+hulEsOKlbtlfojWL0q4Er+GB4Z4My+WTt27sX7BYzjfLHL0jlQHTB6vCfYl
qDNbBaO+2YLRIGD6EJx1293s8ntwA5JvvbLj4xoELb7qkxUM+IWMUIgbGKkqSdpkzSSSrU32mfXE
eR4hNV+Cczh9eFI+WsjdV1aBHj/o3c7asXh/1wvZ/PuUtiEafbpooHYFpORsqL2DP6w4kI6hvNdo
WyPxV552QKNtAnWvU/6YcIK6ay93+MYB7XbnQLZOoCRGUUFq8vR273s7HUo9XOvHzJpKaoHE0d0M
WcJRM58/farmCoq3GBztxZ3v+c8cq8INY5yHR+eahw4fMz6UyRM+3Nb63tgpjFT1qUjCJ49iIfTr
5X1tAR2GIS/EtLkryP17nS+gDeGm+YlP0WDFYCcL2l3SCi1PSdU4YHOTxowIXsFP2imn14j7Z99U
DI/rH5u2PdqPVxrxPCPktQork6V8N0DzncET8thol7epBZrNsx6RHdt96xjDgUXVDC95bGgu1cDy
A6AtgNBXY1SFrv2u/cJzS6bYPlr0MDCRbdgO6ZZrct1z0SJ/qIyAaj5WULhBecrtcF0BNHKdu9X1
dR2sgcMR4dZ+tWGzNUDbLtsbPHUV5L9uemwzoJJyZ1zgruhHLnsaGaeMH1tPqjF/mXrtiabjTHif
rUuGBJOLi4jrS1r6nn83r4W48c2SLE2JAY1/lizkvpSqoyVFnhwk39T/1GXU/8cRxYtSt5WGT41n
kv6LzJY+w5MlkZxVDi688k7gqb2bo2oQ10PTOUkq4Z7kScQ/8UX16Weq2pBPKLYjSOO364hGemEs
LAyrzN/3tNfyn5w63ePxHBDxbFpZzjIxmg0iDQf9Xbx0vO0la9TruC8gShm3HYHSHF6CjmNX0DCI
eUWXD4J18/v0hbvWaxzIyV7KpuKVZehZ3uRSF4McQbH3kfH4AOzdWpxQXhOWQEAVa0uzKWGWucTu
4adXKXgeEC2wW/+e0gJISl1cf5L3dAwVjzxvtSRSNpq2CZ5Qo918B/o8SjCh+edSjUgg2SCce30I
4GJaPzZ9LKyGjnz0K4/+0Bahr3XFTHsikrOSgh6MFwgn3lV28mqZYMXSvOjdZu6PsJKH7wBn32Dn
+LdelqkQzRU41lEgJonD+qEOPuyts4NHM/BmiXw/t6PK0q3EIU9TibMxcvp4030ra0YLSIItqB0B
rkjFCpLNU02DgVVGqeZATiQUypETngCF3gmC+cSO9uJaex5+37IxmrOYStEs5mcoz+IKUfaR2IUY
UM0vdGEWGxIRRC/26WXR0QjKLhP9PsKxCmza7VMX7b1YwrdahQgoobWp11I6L6urjrzeikjALYZb
8dx3ZK0TSYP33FZLYdON6ELTLSXGEO+eFPwTSY8SJEau5fZwHqv3VexOldUwjnz2wV/t8gsv7E5l
cBxdHLe3pnzVgx3BuxyBMatEuvjh6mo0BS65VmFFhXOPEDRvJJmnYCQI0ILk6kyGKGv8XjIG6YtJ
ebW99kIj02IukBPB0WhYVRlQapZKzI+e/Rzb9k3Q9sxM4fbilS1FJAy+mvpmUPnzR9D3UcGYxOaS
5mB99+nvbEeysLGA5aN8FhE9S5juGmAShv+8ZRAbiE6QfaURf9pV69mkyPPTPNaUMQn98KbxrPYX
hwms6kjoQD1aCrpRQbZjf37zO5t4KPqejiV4ihe5uMEEEVEyk+EVKNhrFSJg4cfyDgpeJuXXcAPP
tcuPcgFozMS6OjWKqOwwGAVrDJ9GjKFmi2Rmp5uXE7JmW2raNAaB3fhX1pE9PW72mhX3/GTAjTxs
TN6TUIFvGYZUMQNVm6qW72NzoL46muQFhhvFYwd59zv4sGZ2aeaNzpnIXkkgUxrMLxK6LmjiAn+0
ze2SOJ7hMTwOAE22+faANRbG6dhZjPvobscbIqNFMs68iEk82tLT8gavhqU3xgEmUfHSzxjr3OKw
EmPCIvZeAqHok6xoRleQR5QVo8eeI6Bte5R2nwpuXZb4QRVYiNAjk4sL+yfH9PE7OGVHjyCiJQDG
sEO/dNhsGzjAhffaBdSiQcHKS+4Bq4gC7u46Vz30OB8KFpSn56SlPnW9YVeaapY641nqhp5IWzhv
db3LYAtOivzB1UwbJYWN22kui6RY/WbJoDUgzZVu62VOXozaRMysDaJy2GMSaUeoSjxA19goSJuf
fjFy8JNAph9BxyIGab6q3uHAX5nhvcV3f5nf+u8PMXZkPGAmqhORP5qAS926y4fNGlOMJVBkHHB4
oxmncxrWHKo2Hgm6iBoQrWZBgzd6ywoUZGh9n6K38/5D/zMsF0R0bg49S7hh81/mKyna8/uLmepD
mdTaIYtjvmj5OGButnpJnFcy0tJQPdchc1yO5zYNNuaOnu6s3ylB6ku7mMwCoe2MA3d/pVVOc5qz
Lm6GdSoF1zBEaIhUNFzMsXzoilAf+x4VwZblK/NSUxB4BN0aON5oNgbQEau32vGJz8MG2O87KZfV
67GSZqo0BTOIYinecZZDjWRxECTuavafSmlzmGJ6CC8GkNf7bkRJbAcAGbB3SYxrsifUcvN0JNSn
1FcWDTVizp3xpxxRHNwhh18Oi0SVIUaS3pFvgYpQ4wmp0XhIPaCRYvU2L8LxSGll/9i0bc/IBfQF
tIeaBiJ+ZHQJHDVE0cbVspbBYXgQSY7UevQ53qLr9WTzWroSEwDwnRG8DTx4mb31n94LL82AgqbI
rrMFVghLJRsM88E15xp2p5mCTYgBDro2asClEdRlT7+OJX88GYB/4qkoOSSQpSWGQbht4Ntzin0Q
fECOypVObr5S/vqTMueVRwd5uwPUhaNVjY2qjOPJK74KiDrcM/wb3J8fEjNkAwEIeazIGVj7YL1g
08JZBuNFwrmLVXvkf3mI629Bf1/IbZ98h2m3DKCg28pByQEc6UO31zLx4XZyI5s/DV6RZTsI4z2R
LONRkeXQlzHqvfZyZkobig+G+ZdnTM4XkzZmOSXKzTGj4/UW4575YkKUIFAYggDYpGR+UbjFEztl
Yf+6wff93BD+mVztOIJTviNgfPjw93s7Yt8ZdaL1hb8lq8Sho/wGOYnRwMHkfxVTyXuSspvjqJXS
PjomFUyEq8VF1TC9mJgFo9HwigBdNJ33UMUT7x0CvIYYl4xNbi1IqpsTgv04wBf9h4OEdRPP7R7q
Nroe3kBwXRzNCeUCh1dbaHz4sD6v1/++ncvxCE8KSSA3CJ+Twq9KoTEEAj1eUAoJjV5FhA2Xb6AA
mKVXOI+N223juAPOQpDgMOuBWowJYFZHcVfLdmJDApgTlpTNmD2zWR5Zb7WvDGD3jZYFZJzKXAAv
s2RMn63iPoRTzd2iWvm8z1YIHRL4fAvMn3vy+69sMK2ZY4JZDFT3VUoAeXkHlhJ2yY0J9Q5Xrwz9
enmICb1Xw+aGQAkb9R/ENEbA2cVudluNpzb7IZrdsUffvWnwdfqJREPtUh87vvNdofFAbCM+ConZ
GNmMjqclEvKzvaJc2Fw0LT2KP9RcslrLsB+O08GCPZf1KSWyf+mrzpSkp9fwDM5wT1w7udMT0DA8
pf4tcliijTwaRTKFVFT/ta63WSCs+NEiKpfwTMMIc4QMpqsoYIISNXF16sKAQtUj79PI7AhC7v90
yqVSsKYSNgH4MZrO0pOMMYZ57XqUScD7OJgEFepzfN83JGqudao0AmgtUX10uj/xEBcPzC9beWhV
7hHPoAywehj2UGWw42uBvHKcCE2svev9cFMKxF9nXdGNavFqutaqxt/TDwBBbZpWSrg7pqD3eKZl
iwUwV91XexTnNOUyhHXaKNRtByuaTJVjMSeD3s9c2ZmcCKy7b68dZIlvSvpbgXXIOzZ+My0od575
TRNpvspLoL4UYfPTB0iDM93U7Ydrk4IG8L5XuhGqsqN2wO5hxBvUw9D1YqdR5oucTjMbchHfUNoI
+10Qg/9w+6PBlCEXEr0S14AeZq9wnUkUMMGB89kke4PSoLdRZG90QBGD1LAT10METRFeEVePHYGc
nammcEnGdIoxNz4mx6h0wgIUZNIqD13qN+OezxHUuSUv9TAzh1eXzG9mpBDYoaB/2cNGEChjBn+n
HKFQxo6+t1Js2ERbDvB+LHdzFkvlBsmx+ZrmGlvZ9czyV6Pt7v5H3HiBNfqDKxk1hk13Q9ipzcwI
huGX9tTppOeMhJHkiDyo11LeMr/jzxsXaId/eGKURn5spAgFZUzyCp7d2hE1igkladRr2nxvjDUl
YGGJk3hkgKsEmuqbSgESd0qbEFJp2w+lfpzDkvwZBRn91JRUarc+80tpFjwY5vL42zSl4iSzhHgf
AJfO6LQyAxDc6asXs6PLBmqj5DF/bsfugPWq2hMyXwu3CDyr3rzYPBP7hLy3VezYLgbd7+CGCmS3
hD1paNDfMlbcfZru83nuQ5wi93GJ3p5AUGQo6lnKFSy8PTqG8TRA+x5yWPBbwhxEVY+GDEK07vuo
VBzPFIeacXnlPhlak7q4yNwIzMW7g8tGbsckyEqjlZ5r5b+ATvCOnKYScDP6vq9H+iaooZmGRVF0
K9gbSg1zoFsMImH0XQR6jxejbFtTSmNtCaPi97SLEa4BP7zCOka+qoacx+dAh57Ae9bLX63LJlwz
3KimU65/SDwHtNx2/nM7HbvVhXXzsISKbJsoLlMteM47V240me8sNuxNZpyYXomZSuyszs0yEWIm
34bLcznjIQjkR+12MIYCCsKolK2oz4hFa+FGxQnQqkSHjsVUewte8brXGTuQdX00MQb81el/cWGI
gzQDg5flQwVYZwGv9TkBrtfahLMMlptkALsJqsgti3y1BrPajdeKvHiveCEuZs6EhkweDkaaXORQ
0O0U6HTuev6rUpniqf3G0re6esSvpV4nsEFJ0xSSh/bLNnWJuzZYjV4Itr23J2LMntDgGssVUHD6
9tKXKN+ml+gLmhgv3/8ETQ5Z7NcJwarreURLp0tPtXD7tuJgWTTgqflvpRTsgz4o2n4SZCftthEw
fPg4vgQwnKEOoAiw4WpMd3qWgU8ntOW3FodubpZhpUufRN1meRXJwNTshTK/1NoY4GVrwoqGvMxD
paJHqN12NjCQMNvhzmbzkt8JVax2vWYR5G3EgN9wv3NkDR1l5aPxTZ5Ww7QILYXupBPp88O2LeSi
on6LY4fykPTNq7+tFWLbUNMs5a4jFsONwByq6w4d6kRrWF2k5Vhyffz8BLszd8lmfdAqDGEDWpfW
YRCzOC60NqVpVWzwiMA/1ENrsdHjGTMA+Kg2fCyoaWp999ID2oucUUVOxR7GQbbKYeLo5JTDwNEl
Kimbr970uahy9JF4hIxD0oM1a7JB49kl1UaKQo1kJghrH0MrjiA7v9PM9rpBdEI4bTdsmB3Q4d/t
jL/shjjd1jO6aJBruDxwCrUTlXZ0Tq5GartwvuRoTAuOyDS4wfjRROaukEQBCBFoo+7DzyEsahXw
IvbBEJmyrSvV0nHgvZBrStPOvKuYfXYxiqIwLMMYWjmhr0mlLi21fUwplN/vm1F00rbrd4hWceRy
Cz7Rvyiv/Bba8hfwGiYre8/YV/3wi79SwMz6MBBIbUdEUF7cZP8ZaxeXlO8uzjFXnc8yQWsebu80
qXFCvnulOl0ekUmfpkoRNrA9e9hSL5tqjtuxEOd9k/Txff4zN1VMPhyD0jOhsPexQUVdype0H60B
54BcZzrpOLRvOF+oofsERzQVq/tY1Y0d77miY+p6c1vIQhRKoki3LZF9rYCN0FV65nqtQ97dYYjL
C/ODJI6ta7JlG4ANS3JmiQ+tmtZbqXpJDtUOXfOq5d+maHXJsUQGCRxpzAGqNs9PgmfX+bHpHFU3
vU7IsCp3RM4HIW52204s2iCDKb0qipyfCqlGafv/8ml7muT1Tp7XqcRR4ewhVob9HUvsCoN2MAyX
Zfkqcv7zLRmBkPQBoq08p+azYiYWk7lhQi4SjTg2DnLW1GHqc/hy32BwYftt3J5W1RTL4uXvmu+F
aVS5qv43WpQ6G9z4GOXioFXJm2mM4yTiu57OPO9C4HSTGiq29/RqTcWgM5m5Xpwk7LSMw1iwOJCo
9Zj++FyFRAmnj9yo5LOIGuandnEMgJbKbZIAeMy0gKI/Hs/f8eURqsGFe2AvUVA4O7deDQWWnYtv
Z6LURa10JGwnAOtivYUQUtuXC3pZBOhFp5IrhyDWbL7eiBlMl/pV/Q8HJpROxbewyd+iUHcqihE2
LG/uCB76MQryum7DP53D10lWDKcRyhL18J0HbTuunPFNLubkaQTDZv12DB1HOYUdvlsgywjYtaF/
IhzUGVRQk0xnhnXDk83UzDNNTpfvzUyCFivyfcbVeEUY0LIGN0VExQ2Va7uGJMRKH+ccEPxHutIl
ADoYQjKGzqVPDF9sV43GkvdLnXmHaUu1+2o5LnBvf6bl6r24IXIGfp7vSnpKlgzelVmD5iF42oCy
rjwMTABMZznVRFHhp3lQodgsys3/uQgtkJAdTmCU8d+T8xUnfBH9WG12rFZRxhbXK7RRwBwpztYQ
PlxolNO99D9+4zOygZ/GqLxvN9nAXUpiEVSzBJj+dxTZ9/2cyMybOjng+xw3ryDFaVuSXH6zUepL
6WbY231Cpf8+kyYd3gdp7meNiGIbgv2m2lmmnKFD7A1jtgfcOmhMncgOk/ern9QT3iKaluWLM4ZN
HTbJvWX6hIYEQ3NDfmVv4NU6CfP5PjiAfZGyKU7N4NU29OjNZd9Hb3W2fB9zcdF2hA963UfSdFbL
vHcp0mqtu1BhzrsqSfuyPvkr+VeKunV+1/rOC5V458Y88qRuwX9WLfUmEAW9UGcgPHM356kCG0Gy
XpFGUbVGFP3zvU5xKiqCv12tKOoEQRAfiXVnUHudwkVYoxtKjxoGe9n24aejw001ortdAZaoiP/F
EIhH5zZi9eSlilQtXvlV5fMkQytexfvmlmUlly7dmIJ8bmeCMTapfNCvDZgFVfYbxL+XRk+brXLU
yJuXQiUx/MbVaXCjnHfkWIqVfQgWqLrOBXujIJuK2aKPLMoPduzjWWDl6cqEp+QOxmxa7/85Hovu
mDI0+3HaonNfAzdtaSHacn/xyuBrK2/rjnNqBaZJlfIHvrOhscgBFVozvqtfmM4EQ81j7+XvkPLk
+y6gY2RGAh2CjAVFdngi40ripoDc3uc9mWxmUhCgt1AA7A3CzvbOB802I6rDONjjIVD86nLd7p9h
UrVoXlmmKopUc1MiVvhXZHoeLl3T5s+N6yw/MXVZuKz4oE1h6qwWmLxkauaL0aMMvV9VCoy7bVfA
oliLRKI+Wd0IZChLOmOTKKm2Bzf06qgfYDy/BCgEPmoIb5YIOPCHFKknZqc3I8ccXhCZryUmYUVc
3PW7wSKsRp/b6LVkB0Fglpreb+xzOpUIsUBv75JrJY692tiNbQBzuOcbIIJ9f2F7vv87QGbyK3sN
HVLQNbCJR0f0SgyHhW5mwvVt21zi86fLcGgVBUrkr7rrF+Sg/QirEVx1zK+Om9Tz8CUjHHjCV0CB
GzOw55KF7JD+61hsEC005RllWUfh1UGSeAP1hfXRtwp98ypwMTPAUOu+yqDZIeGJS6BMVQ+YIhtJ
FYtXNnhwNwzbnt2Mu2yYoprKxvaIkszRkQ4+j9bAgx6NowOxRjLjh4YqGDJhsaGFik8buEMyjhnV
S2MDo4oZulurVvS9C6mbkW11h9R4b6mfV/0w/Ku7IY8DmrlPStUcxCUNzQv8U69MlBwQ6vawZzRs
2kCRo/f62vDdPDVvAyxuIUh1qyhXTbkhsYb+gVFFPdZ7+s0h8hmMahOrQaKhXI06/uE9pWbMwUn7
VLpr7dGWTkjfgeh+fvW7/XlM46osZ3UQ+8pZKezrbtR4zZX3KfgP9BoJeZzVV/LdydOFQWp0z0hd
5m9J0i+7sh0iGLLdsQxgMgpX8aQw7UBzgz00yXpwy1cER5ln+nCMhcEz81P2e05PPSekdf58iAWE
oXWvLSXni1jjzx6p5MxkzZcPrlt8mRITF99pZZPGxCZvW6GX3WeBNTvWtfdE5ApNoys4HN9vAE/9
SPWuz3QTsHedMT38St69+woZwvchgx0xkch4BJOWIjdvQPLuR3fu8jWJdJB1rtNDowzNjmXIS70L
KTumoCkazJ+5ParflNFU3blkAqifibgy4ia9p1CEOwGhDmuNlzyHGgznSaWSxuwyjkx3lN6O1iQW
dltgdyPQhEfxE1m2GntrMnDQdgPd2xw4llGUWM9qbQmt4YZT2l2DKhawa/z8hGY3fODgUg/pZJTs
8cOk6Sa95jhBMmTZBuiXJWF9t53lO9nOTlO2TzujvIl3HZVB0zJu5LLbrGuYFFD06UwDY/o1/Qfh
pKNaPVIhkUMHvatrnUkDC30slYFNcJpSABUmzrIfv7rkSCHp0aYWPwKBjOXfgRsqGCpz1Cz/nPuC
bqh0zCedFTIYZX6GrZGfyXHV8iMF2vEnz2Z0vZe8KTSOAy/i1QoCIrHt4uw7zdAyKko1TXFxUMTs
M0WUqAaPrge5Hsb8NUC3JChS9llR+7r9685kgBh2yP28UcuixcqAeMGO+J3Qva+SIVVOXtUzXkxh
35a3HQL6n4gx7Nhh2hcCNDlbQoLuqLioYBtRL7pgxqHiceQMDNNr9noipClo1beYAmBIDxW0L5yM
DOlI2XXSquvgmDjBTbn8aJD0APp90fxQORFMvZYCAUHmfGzJ8eCMBifdB5Wd0MkNCuITy6mynfsG
Vt14HgKnnsRmPw+sqrWW9KIHjhPh1qahOFmmhZJ4dsiW/37Cc1ekbLHa8P4LY9F34cWs0Wa6/SrA
snF9nmnrjMfqmxz8sDXiZ7sUyVP8JRyQRnibkRJquQqa48o6Es7boo3+/A4W2VGiTyg8rcnDzjdx
ZrBt+3PljEslvstnZ/BHfpbazmDJYy3WDDTKat4u4PA3+cQcbzohc+FdwnMwGU2rAMF8wlG0I7Aa
pe82KdEt/LEuMe7hhXNTX8vga+88I2JZWkMlC+W2h561hoIurCRatFicKDMBBNpNWHoCpo91mGcG
BFdEZ56fYWrhMyRoq6lXAMySRzzRG7dMWNYeKGk3o6TC5vVwu8uUGSCvAhkG5GEjcPvspUyxbyrY
Ura3bPi2e0U9/lvNM8rws7K3xQq0f2U8a1Z44D07fWcIk9wg5QDDtm/QNEzZDvh8JCnQiD9ipsbu
BGgN0MggXoFWX8CM5km1dVGOSOkONwzAfCIzP6uZOJpHj11GTIBmRKDyPr3io8RJz4cKKBgLwrdw
ybaxUp7dcVQ16v0PkXgHiatIyPT0S4Loy5zs3CPcqrElWnoM/yQdl2xx2icOf+7vR0irUuKRdGmI
6Rf4nuuOzPBe/6BYC3EbDjEluMISyhBrv9OLJKAv4jeGVGbaccL0WI4+jZZAet377RywNEP8WNg9
duwlSig8ksCsEddNOaKYmC7p3DwrWljO0GM7oceXuAMIQyZD+fHu09uln2ouqODReeZXki6qgTAc
dQwfWtujdPO3PMjDpEF+C7wO7H+MxdwTMHlivIKXqi8DT5+HGmU0lxm6W0kSRJ7MJbzZq+o/N1FE
9NbwejxXTYNCtEO4nOHd9wxv0vd8BvHr3eDr5FW+dupqHt7+/Gvt9cLR6F39ve46STtJF8D2dTEX
QppqzyOA0MlPdIUacuAFsCJDDuKLt547mBaPRUAwjhleDsTXoURzhw3sl5pXVuYZ53F3Ev/gUqZQ
zbIrosIRpYAV/3kA9UjF1U3vAIHW37cT8zaiHfB3v46kvHbZ4Arky6e3H0PvhJMkWwR83Dvuz7P7
DfDvjPEeVLVXskCGzS/1DXJwHZL1jfRPrwjjfNUXazKDeIvQF0JNiKoubdbVdmYpdgB+CDq8GzS2
8bhJOGGz12JcJjwcW3ana8Ezxm3kaOTibPW9WT6ObIDVrReOXbEdFQCPZTWziUONDtOaI0T9hSWl
Vo0gFP1UIQaXI1KPaD/MG2lguhmSBGtMlgNodbbRKCoUtLnbKpuHqAoJsym3TgwBABW9MZOP+TV9
ouTqlnOeZPGhLUoS5GYl2AohTZAK+RvAT7atLKePaso71v7Z0MvPaNq9gh93T0HHEKIqIaBX2v+u
+YqF9z4HFkV4VZdVT1be2fG+XqK/atsmUhnCnWO0ssrGgE6ZkYIlw23Tttt2qSmWLmyuuNsBVdPy
lpvv8KBcXRglfIENI7zJ2JxhSmysnIVWtNXJX7o5W4bWQLYt0f79tcbQ9SazYUcdI2QZrSQt0X1O
wTrZyD+yNdeWDA8C/+GTUUZUp2Se35AP/maMs235uC39/QQX8nqGhcezwulrMsft8fQLV4VqhM1x
PPdGSQJgTbyVQ2HJV6KDO7e0K6pRzrmrHBfG7fRmKJSysz4kVwOwy/QgzajHrRXe0TwZrREPLjTe
6d/uJve68j8FyPt1KiJgKjzL5Ldql3wkMiVaUNRFTdSpSMmBIjTRL06fgZoBHDG/DlfIOZPjERVq
7rmulKI6UHQaSa4VnB2EiYo2lM/Y1I7q4BVVQXE4peYPKRxeAiTXUmRC75LMIHzKiWLaXCtk4poB
xFu70YqUkWiNQvKZruov+fhv7fV+pKRsYwTNgGOpbaUtC2ymuTh5NJiQxl711H6Betf4oMCI3mO8
JDTKtmLzLgyyyCN7S2P3TDdJ55SsG0mGw8Zj0rzOHrVvR5ZnVfcoGx9K788TCQAquBL2fTAgjYvm
571SwwNoebDVkzhMyCMHSUXLvFjmOMjC5ka+3Z0aT3x/hjl4VrtlId6I4Qpi/3h5TMMmcVWK73jC
EeJ4oTpbJylNgGxAxZA+j59ZfWS89xPCpAKxlkobIF8dMwvevP3Xf7dQ52CvOvf08kO/xYXslFkU
Ls1zl4WvoDEnha1hF/wXtUUZPaAmFgOD/sloSnReclckcP1Y2jEAcFhDqYOPvmJUj8TjGGG8txMk
9UWJKOOLsbLBz0WMRmYBFzowusseFGihBxk1NPpFIw2RdK3obrKOlSasB/wko/v88xwwwiprvLvj
mKRrGQJHSFwfnZQMmdtx5mpq1pcetLHpcrWIg8zN+BZNWMtoZHGU9v5FCJGgDtNI+5uVs5U/AS2E
nZVmNGu5PCP36tfo1zy7Wgk0/Id0m1fKD/V7VrQukFa7SGCZo1H+IaJ2crqNSg6e/Bt6sQo3pOqC
ad9klOVFgqM8FqJ9RR0InY/bkV6XE6caSAC2Cm7OUxT2QU02rVJUpVC9ALKscUCeSAw3vec4Syml
PnyAnDQOZUFwaY91rqLckIdEGd/nAl408KskuXje0+RYq820vOF3cEkVotDqXFlIAPZjgC5X6r5V
lUDKO6HvOKGWDlBhOG3u/vcRor8HS+uH5IY2sQ+jI9BZqs4KlkMIPdhVU/7tyshREu7iccvtU/hF
SZrN0aoV9NfT5K7xJ6Q+ToVdgwfH6tA1tzCz2wMFg3zwU6FZXUJBLEdBqRzreYG/k+dNzcohTIKs
flLcxtQXH0I4ApND51qneRuxdxX1hYJPj+WXTGTyP5JPTQi0kg9r8huuOC8pclTAYObIYPE1DmvP
ceTKSD+PimA6lhcWtHiXfh1ghFOWh0sh3Wl0f67/KxBR79GEJFc1aI1SJkVOY86LecM4+2oOEE0l
5ILInisc0aoWnNNT8lNrnlABxizTT9MRPUjndFd6js9ThUrtgYT3bVt1RCcuyvLyyOqWjVrDY9lq
9OmzWKaeLdFeJVnWLcX0E5XbMUmSY/w2nvppf/tAiieVY/wVHP1hnhXjMWqMAQI1Kw+ODcW95DeM
7+bxfk6PMAhvoooe8EJLVMNW6ufyTzWXEikmt4FTUIr566wQVkp1Vs2mwlL2benJPGzo/OGtAWjv
RoIHFsq3H7/Wi1DuEt5rGfw9CRL5UMJjXb0fvksg5qjNqRX4lxIL40jd2z46J2VBfuUTfF6rTIt9
5/fucKmHJ5kYowFwu1PGmPaCauZpg/KHfeBjPUOLLPsLLczaaxzKDoz+C5xvRV6N1hne4TLML2dC
XE/HHwsrzzGG8xRiO62O6iCPdu68IyP7ydK8VPXokbBn0XSsRomDnREOKmzvAMSpvAfhCIC+0Y0A
3calfNnUS2AGphQ4p13BtlEN+Zt2g5qMLAv1UWdx2FKBqKr4Durx8VTeZdf3K54xzzEjriWW5vr1
c61HEIFUcp27i4g3K/88ji4/btUALRRUgaS199qVFaf63bPiHAwZpYDIN7s5VapDKK/PQcJfz3sa
jIHoPV3EqyZzhqaUpa+xWPF4qkJTfcp+HseZ/JIeflnFvbAqCZZm6RdqZEtv0daaUWdY+znSzpww
cvciPMubhJHkMlklbvXrjJr73MshT8TkwNlNylzFsMFR87yOTXYNL43lBoNlz1UREW4fBLZl7KUe
JYEmhwHv15KmwFXXWD8ppvbFl1Zmq6G1daLOCQt0jefP4v6G98idm0n+tr5f8ZPtwcPziJBU/rbK
11iZf2j9QxbPg4e0PloxRls0WvEDiDwGCgbapkA4yP2LhVQj5jwLWmliol26shPFWdmdQgJ3hK+q
VfYHyuQsJx5bgjVkj5LtkpYj9gEFOZv/j3+wu7s/A5zSndjs1FOgUP8HHjL8OQUFM4NK6V3YNqVI
lwjckAXsQdX9ymHB4EkIUck7goDNqPyFJeDCdht6LUWPIUpjadetb83l0NBxsnAN4xi8DZQ8+lWP
Tiogikl7ml055eJU5o0JFbmjcyYOfIzsvMdPbP7+N39MQRQnYPqRnyuyRTUGJS0tvyBrohPAJkks
JPQvFTZSW0A0YfByoqI0EdPq6NQ2mGZGVmaTnFuHCP1FDoUhsWbwkVNHhOb0Sg0arDG25cdzPfK1
pyzQjjlUD8V1N75amhtTJCnHjLABqUognkGAH2F9PF5hPNnknQP3FayUaiXZwPMAcTPdlVGzjlK8
CcTcxkCgi683BLDBvX2XkAwOsucx50QB5h/H1/mkhkd3B8JiMznFrqXRxEp1hXVja+gN6HJO0jjX
fGcv8VxwNvru7+hYHLGKlIvRmDwj1HwPbsEC6po9J+USC5mrez85JNW8FtEu3zpJQ0SjOuQY05Qp
T9Nk5JRupbrfLY9T3HjFQy6BpUP6fJae0wgubozKD9BHSFrAw9xMulygVRT5zvNqg2nHiVAmgiOK
ZVAFfw4kYssUWEOLUFUm2U6urkHW2M7E0PltlxRqYl9l+ylXR6+Ld9wVwNULFDwv7wo/m+1WTUpC
J8llzmQXDSJRwzLwGrk6QRvhqX7gZxqSI7xQoeQenI3FHTzaQxJ7y7zxyJrXkHrZY8rh6HRl+kGV
bLS5dIeTphh7GoEnhtCI8iR2+qCXHEVybzSrvFW5nKsySj7wBS+rOb/vc0eWYeuym/UxdVkG6Ok5
swBxJchY/zV2QsUNRWgM2B8MTGTL4HPxmTFglHSfYphfw7WZ7QZinZ/UNGlolmhSuPBcQ34SDhS5
3hOxIfuQuzs8q8yCNk5cwtCHxdDWbYXHv8Nys59Co7ygUvkR7VFezzQSrbypkYVaJE3dIynP8Qej
Y/NOmeTrm+d6MsSKl0eswP1rZRMiiXoSKnXQ7S6nRTFfbA8VsGA1WeSTTEcQya/F4ePtI/LdpMUy
oIa/HWdhOblNTwT5M6M3oWMYoF6Ktke7HdmcjoyKcGGd+YB5u/65XnBu4DFoZ/VHah6wDg82OyYF
txu3TqWhFKcPl1cRQnRMM5yN+KvDpVZmASIy6Um7b9G6Y8Fx5DeU0CEiSQmXxJhMGpDAZ7i4NC0l
D0hU0p/bw/T0Vgqank8H8d7YV2Qq4oe8EmU+y9vog6rNKO4cYBKR1r7T1qnfv3c0wvm82VHeLAin
LGVAD5OATZ+biEUB/mZtOzLRC8S35AJLbmkP2cBofKlacMAo1AYgyTxkDbXkyivFIA0Yfq1ELCWy
ThfjbWtg3lrfwUxUukG8KvBLFvwGo3VBEUJ6jxR9b7EwOHhA0CLiVqrhIYlMjiV0lcjiwu+0N6g4
thhQiBuSh4yMbYWrhQ+C2LvTx/tkz3iB9D/RzeL5nvGEyWARshnKoXGmVx49b/1eE1+s/KJCFMCV
Ke019pc1Nu6chip7qU5y8mkkcRyB/ffbktYkXogZctXLK6oRfiNPY3WTdfe9qsOuOQRW7lNGT7XM
c0uJAGTXqmuBeL5AVYs9GpiYMNVkLMqykyjzGxeIEnXgZ+l7X2lEFkaWas2zH9hVc6AtW5eVBqjU
pGfYsCheQcd7a8+iFYvwu8AQUdmke+FF/nAIE//I5IN291CGLSooRofXiBloIpjUcVsglr8dWwzA
Ye0b1CiLj51doutRau9KGyxeHi9pR8EH4O7NhiHQv4e+2kvhtlmMF+jVgl8lNFLpDLmbNEXs6Nl8
81PtzMlG1zOB1mYHlbW84pJoG6Ias450VMuxveCyhcQsXkwhtcXiCmJtO+QCMmilpvVHrqeo7jOU
DbdnOoLHnU6/IM9rZWdTb1fVfhGS5m2Vgv30QkUy4IOxK2rpMZhyTnA+XI1/2pzsN/L5tmj5ADPf
/DvtvbDgVVEanlJiYl4+JOzQk/893iON7fS8ftFYl0Au3lp2Bfhw1dW9WYhJig3kAghkzh9/u4Tp
YrYMexR7YUdERsjLKX7J9di9X/aJLg16Vpf1HZBVFGoC/HD1BMyUF7T0FXJC+F/P2eT7tRBmC38A
7VcCD+hBELfGDA3lxfbtf45ln8FCp9eDc1nQTTfcOJpxnjopoyfTko8jYb3o+WWq3V30n72MOhTW
E+MysfJCEGGcpXWziGl/PGAXurMU1MFVQmfjIQW+Zmc+cWR/7JntkpSbACGgsgLDvd1jdiHlV+2k
mi9BiIAOrIWjIt7YAn8rLMPadqk4PmU/vXkTxBnBKfurykmJDzL/58ry0vNOzF8iM4XhsKtWjQdO
yu5A/vPg2UINZc1S882j+xw3dQlGQv+AaohX4hnhvw3J4fwijH8uZB/19rZfF6WxLIDeP7cQsGPH
+TS8bN36cFuuSVdGeizas+aGaK0iuHunnVaMyeuXSsM7Nskn9mXaAR1+EnOycO2qGo1+aaiuo/Ym
QhVPhtoyaq2asX0lXNlWNeI3lCxN2iPu2IhVkfbTE8peh7MdvtxY3YdGfhL1qsY6PHRnvFz0fv2S
ILbBPk4vVLZnIhcFfg2fDAfzTF5J0o/ks39QNSbKh0m7bftAeDlu1Re1TKYdDcMCh6gSDvuzkaiR
kC2buupbkrSDE78qTGJ0giGLCGhIv66y7BRErokV6ITGMEiHoaLK28G34heFFGGxmWFHaflLWqPR
eNHAX7iY1Nm3SzjXex+VJwDaajF0cEHd+/dlPD4k8xqazTkzDOzJHX6mEgOrknx1m7XOZEy6TSxh
+MqLEko9Wi6cdaT1SflSRil8e7JLZwGJM9yat1+PKBaARa8H5wXJENBWmypLDWo0/xxBf7D5BNio
SWvinp4nwuEmvt1ysJPUx+QKPkEFcNOO+Kazv2EdUJMZLHYIEpaTlGJ7bpkVWbH3hfp1mmHExF0C
ICWX3reTYqVp5c5TwMUbFeZXgfbOTMB7bkvxDsValJIiL0zZnVLlrLg1L6XAx6fi3pWwNl7qqGbN
ERi60ejytgmT6NWOmdRZd6CGGxiHegaOqMFoqqFgeVbUaC9gfogar9D3BVYQA1/c/9uB3vWA+Ube
Ga67z12MuHFl2Vltq4MTEiLnoHitdSGPT2FfvaEVy3ZS0gPQafN6D2FEwb5eUb0/hEh+9SJdeOX/
GVbCq9f+JiWpPpNqMm37XOo8lCvMd8r4aBrUXJD0QYpSr77sHsJfl4OiLpT0JrLw0i++WrAgfZNe
xKyoa8IyRx0WOiBNaDMLWmvEAKly2RlmUMvTgMlNbD8/6XWILKym2vFbzhImcsJN9IahGOCJdm/X
2zRbWqv6TLqwAiBYVPbAYEWJ/lrMFU8F5iW2Jb+pxaFMcMyz3LDoYZsUPboI+OIlPLm30N+YsBFK
7osaDs4aglabHBmdTb8ZEZUmjdvJGxgI5zJARxyXLkqtro1qECeO3xTpHZ6PSNKjZRmFeIJontgG
Wzjx/4QPcA0J2+BgAbjCjgAm5UUvhvdjPpXPmR8UO+uQh1w+ovoOT9G98GzjTb9pjbq8EQ2ntvRq
FSQdQOE4bGfJ/7e+X1DyC/kPNkBHJ0mwR6ODPmiDfEz1AmTTlCtdgELWMlDvMk+94P/T/LVt8UQi
lC2dDTwKjp29Phr/vqCoS3M6Ch4KUDVKXhFnDK7bTQsEhU3nDRExjfK124OUmITcWNGJzXzX/52i
HQk+OXhOQkMVrwmnDkSQDAc6DwEl3VbEuSBN6NEaxmWw7Tao/h4Oxo/xm1iz7nt6caJgBKDrv/79
dUzNUY/yj9gQ4ikmX8yyWgLlW8gxyhEvjfIehkPB4dzofyECYxUWWhQCOSFrAR0wEIln5IRbutrq
ZsaWLWcjoci7hsi5JOs1RqVJfJGh54raVAZ4KPfWGQpwJDW7dNQ7W1cdd2jYVQoiTcVyvje0/Y+v
bQ3bJ5UmY+7MFjqDTRg+el3Y9C+XG1uHESge0IsXcYh8DWGkjgjt9/xGJc/z8HzqkZ3u6OzKFuHu
GScS9lrNjzoHNJhMGSKdj3K19iMUxcKmcXETZShDX62AxGXvaze8ngmkEhWMiLH+jP6XLNO3LoLx
Ti/E8THIPwwiBfqChqgSM8i2CQ0pdMYlX29+GYNUALz/bpij1fs35/YDY6RzQFxx7tSUBAveYnIW
GBZhIKekOTyN/4FlnS/GPLFJ0xMDwk3kvaSM2Kd+3U6d0MTtvoZbnYG8nbudaWs2qF0+xZJjKIBw
dKCKfKZg2f3DmWO5JcZHmOpXfMqlLAuJKT2vXBzlqe05vBFgwHKhyzHDK06/GuIfdRYNtzWxebU3
vTAPtlH0U5YLRQb7JGrD8A90ZxiHDtpxi2FiZWsn66Sc3SGO7CjZxLGT/SzeMVn0GsIIzsrdzHAv
JJHnCPTYqqrQ0VjB7akrNBdN1Mhwn5IP/Flzfu1Wh1NfLphNx0MuEOPmx++awG3JwsOEcObZInJX
DvnsAwjuext0cWuyj/1T7gW7bLGvB/Keq+9zWLGh9qvDY8/sePMXSKIOZG8LjskDVCNol1m8H/YY
onYQ5lHi4tFGjNuWMy/PwSBL3hO0GMNQTHap1XrEtSzdkBeT5Re1usmEbvy+FjxthMBLfyWZgYqi
CTF+gnVCjySWLonh2J7LZytbWOkFEcMzY3ZQ+APOoblx+gEwYw+/rVlNL/VGz6L0rCclPgLSdZg+
+wQHs/uqW2gkMXyQDgDtQHeWgdNOWx9lDrL/MtG/Ur1JwB8prYx1DFl/NrilZ6oNF1Xyohd1shLG
6mKZqAwq3vqOzlrWXCDOQondZu72ic+DvYNYRDQtvYDfn037P9SwlXFeUuGyDCnR12TkBi4qSQYS
4yDyYDSORWgdc189Ls5dVtWcIbcmNjkZ1w29yj65XUZyVlUhqAF+tv8WrT0nVMH3IxJMQbvgiC4j
gx233i+1gwOVWr+FGoAhMDELkABb1XnxZcdlGU+5vaxg2T/P8kIesRYw24js8qIWf/03NBV/JW9g
NFBuaeoMh7dHCOxX33KEYNPcFLxJLYXcDAgKv+94bTmyipnXPTJK/0JuNo5sdkToL0Z5ber6u0yz
TQy6qif1INfDi6+4zeZqwaVZgjdzOWo8mWQP3sZKXLxYoJAb5jmuh4L4kKqOB8PhhB+IfOgWdaLR
cEyLlEVpZYQNtJzsUHVAjFq1YFHEQtwNNk4T2/EA3DmGcPdcUeYrHSW78kKBno21OE37XSlCmu8b
3F21JDBFMNMaNLiDzfvp4t3ZVTBLFLbaJG6vgjXZIgavyxTeZCeICdTnsxg+mD/z4XGvlYCE44HM
NlftM21BM0WstFJWwmBEvxwx3fPo/XP0ybSmd1TUbj1j2E+CHxZqaG/bccLzdaTScoARAI5QagrO
v97lCceiFCjJZgj85h88C/eGK2cL5EVE7LsapVn3ezYTuidfqYUKAQASc9hu3RMxkda2bxtXg9vO
0vRkaEIHTJpXgmtfKfTms7QyqqQTFO7OShzEXOejt+rmI36wSkdmnilivooMcxo6mCPS73e69fVn
Mu+GrxlC83rlnKMN9ViUTiw1LsraEISwBpb0DnQTyElE0Z05lSssQr5fhbA5vif9deWQi4gdh6HR
awgjTxM6vjvT4fwNQQjIoTgyBMV7RIYt7Zqm2IAhnZo+RdNoZ/akruCZl8wIxTh/XfzAivDoDrNe
A728UbMH4yBoFbX0RLhLchQYGYhotDlWO8xV/s2B9PtSeog4rz7Ux0UqxwyYm/SQ8Ib5pka2jGsG
MT9su/GdcIKVtY6t97i9I7u9xOykClIVQwQ2t2gwdu2SfbwgSDpSBZFDis+Sor6EpQs1sbIkHb4W
9f+TA1QQ4BRWWQmUv741MPwysRUPQoA3T2BTymH33JEdkOCOgYVd9vLhEVAc+SbMtEKA4d7vcRSO
uWNHH5dM7nARMTZhT0yJHowo1XDSClWwJE3Bl2uTwXsPf2XPnn1lq4tVKUmeGTuETEe7/xg5H1R8
ombpdEHxefemjTcAmyDc9arJFuF0SLFTr2vQqwkyDGyhafSFjxQ18BOz4l1JaNuH+4AiGPeWt5hl
473hLPABG2Wr2g4o2dmxxNIpPR0J4D33x+TE/aKmftZbzhy8W/NOr+xxPT2tLB1wFXPSFUwGDshi
GgqTGZ1fKsr5PbN5E0Scfu0gN7D2Jtz7+KvuRyaqx2hDLFl7SKYJw3qBRLdUFxoXfahr68JJd8U7
KzguFe+0d/NHgjpdgQDR+j6SCREQCaJL29ljWZwJRFPO7jP04gkO9ASi5Eiz5PNV5CjGKGYF8zf+
K85NZNVwe0EQEJNFHzMxN1PS/FNUn936CgyB3g5Kmy9BpwvgRxhd+uEVHHLaK7I4F5hSY18bFohU
fVaPVOGKwof0vrjs+wPrA9M6ngi4btUCp6o2SnL5o3jd5m3xIufRPdnUtFT5TJ1odk1Izjddonym
+AppNIBm1BAnxevjET9Z9MoCSJEmHJZEQGIKnHIftjx8N9MsbgBfDUE4A9NjSfbHuxjvHXpjR4gY
HtsQWDEKq804YY8W8zReZGwIK+x3uX0cw5+eJfLvqrLGKHZoGz5qwzP9T3rI0GDz48hXuZoWtTjT
DKYB7LPpQDqNpQJAlwJAo26Eg5jAZVxH8RXp9gE3GkYUuQG5Q+sNxIzW94vleohjvyweM11glTH6
7PPEC3gAqbS23MNk9vWMqCZZA9KaKoST7YWrExYmjihU5XzgevNiVz+w2hp5prwlM+zQbFSQNRey
L+V5lqAJkjO0d8uY3DUA00Rx29FDWdzgzJw4UHo2urv6+ndGwzbxoksB4xup3DAEVnHxeD78f7VG
48mg95cYUGTPJJGxIiR4K9cBzK6mwCdJEXEXqXA3idBy73nPqcOEPupR74rkbSfMunVukNzgnqkH
D0BOwBevWMr2BcA+FrLz5a+1Mxs50pz/h1GjH3odm9qHrEmqewnoI+0rhuHII78bdT8Ym0wo4gQ0
jhgEpGvJ0gvmT1Y1C8KiDWTIdo1JfU7i9nPfFO4GkjiP3+QYpCWBxu3Kj0dy/zzjGAsmIFflBW5O
R19k5FK8EqHmDacI/CDdzH3YL3MR9skjiXiYL0lo+PW0lHk0Ieu3fMc+6KXcVhleuyVAN2QMXx7w
P0wwFDKGFrdm3ylLW8BYX/reTSCTbso/3YRpjI9E8uOL7n2HWc5u6jH9+8limmHsp7tW0JZ9dcYv
SwDoWpC7ZwkzgLoOSEsIrX/+OBwpS1A52ORUb7vxIt0ashQwQS6Twv8qUuUgJxpIEDQ+/M1Uhqeg
pOJolpnUFrjA93XeFvRL2bLEnyumqoKzQ3KKiVA2aTqvmkSYvZc9tlDLqspG2hU8TyQ95Up4W776
4GmfFfl2vbGIgiew7LfgPVjJTJCVBZPwVA9daFMx85xaxnMb0Ls8LG4fWr7QPA/qM2xagm/XqJyG
aDlt+ZWOKfNjxs1MHh1mJP4ttwm4LLirffpn7cx8nmpSM/7miV0rjX83hw6UBAAgFpFzi7wwhnlm
8ZKYYhSINu9t0f53fUr9ykfh0ApZTkgiLxH9VnP4wMT7s37CVXCDIoYUQOTr+SaH6FRxNzVkpghP
NycSy+eB3eDw9wHnGo+1vdxpfEmwnDB76QOE5aQqJlaDctEUUTLRD9RPFGyri2LVIhc2p/6wNaTX
KYaGisXXRua9+CUIMFkg+TUeiXNH2bKBdrBjqpjlgATFWYwUZ55DQ0O/iXDRzvKWKHA+RgTPxQBI
+twpG4kBNr8Wijbyg4U5zTg9BKxRKny7081V+XRnUKwdUWxHJrHaVxaKxT9iAY84jMTyMtRn9fPF
9j28TleAzdMIB+R4xMNpHd/jgDEkG9HIJLWTUB3RalItuq4FzWqHpC7mT8zEsMvA+mN7MiBZFeuf
S13gF+om/0cvytkzBAY6Tp4mmKlP/0/+Q6oGothk0fAqptaZ9YMnurPasF3CDtX7NlIzwfyGjALV
Qk61EupUaWf+bJcOyNJWeK+5v644APG5CLKPeAwyKiV/HLZf4hH13f2l1oW59EGlY+Mk2/I4iywS
JJTMiQr1Vh8RgsZgyJRQBbAo81V0CAPz4FOKbUQKFP74OpPLR/wXATHNjeLMybJ6c0NvZMvFFg+n
CxcjdB0xBJyRBjksT2I6oTUt8iEyloEmCei/4rVsOI5XfaIAqJmuOVotSj27IsphAGDkZzG+VR2L
h9e51IQwNs96nyy1ktFT7NeNdkpzGs3sI+oB4SVifopvidA0VxgqNGNsJrWHVPXN+CZC8xdio2/T
jF4hRd8Fr+IM8AZyfI+qoWVCPgyLsPyHJrplQaSrnghzEL/CMQSsUmLuamgqASWXO1ZMPDo6bfnG
7gkxciEBy9oSTupZKmh3IlFgnj4sCtUYadgcQuM07Yrye8Wn/pEPgCBienZVEMUX1NZmJfAteITX
YWfmRG5S4cj4cOXBsUgfQLce9NzTMgHLQbS0IaJQ0AQF3/OF8+eLLKl8iKKsbfcND15PkF6b8a81
d6R7Js0741NFBhkI8h7nWA10wm1nAaO8p31FiPcRaPWwEN89j7SKocPsIK2hxcv8U94gXSmFysyd
yiDzy+FtrtWxa9oa66Dom0NHawOfzdPp68D+aaluFiHSwUldfnJ6ZMlN/p9tW9bL7Nm6fvPc1IxZ
cnjBX+0UKuH+W3CzBPSnDd+dWhJuooydPYtc8om1ZnnXWEHvkLdIzlW58ECBDBKn0ibJE0hIYZb/
QiIcvcekQrALY35q7ap5DoQHzuWBLOrERrZIULlpGSzpbZyWP6P3H2cUezN3sOBss38q02OUz/Il
UQAD4lt7XXegnkYeMhmdD8B1pE7YA1qRNWrqi7glA1MhIcywMpP7Y5h3KjYniPVe7y7HusgxfLYR
7R41aOMAug7ZJQ+c8NmPvrBz4ZkEeOIQRLMiwrmqemXMBEYZajCcgJV+o91doZZdwbfQu4FL8zYL
nHNtNmW9S3ay7JeMcD4SCe0yhl1V0k+GvoUAuZIqEfrpb7QgY9IjhSIlLwZlAbRGMsxmv4su8Zg6
WCTwBHNheLjW6aF/RrfCApD/1zNkLEOyYkLI/6shpZ+qWsIFv4mZMuau55hpDQZL/xu850GSKkKj
l/7bFp8HbDWKMg15jCnIZycb70kRnpOe05cr0whiwFu+xE1+4AQ+HlNRqLbETxC8q8FIcqLN0twE
i1UpkuaJiqU4D1aAbrFBAFmSgho0bovrnDky7M4t2ZEm3IfhLMM3PuFEkhfIa2wrEhLuYay6aea5
D4HrCIqeLeL74L4p2C8ZmAOYM5ZCKl43FlGS2cajWCnFdR3yGQSdoinWBwyJbLJOillXKacLibIt
f7C2JLMFas/vi0JP7vEGmD1Cmx6tUl2P+G40Wcj8E7AiRMDL5w6BcNWYy3/TmmGTMpVFBaJ16Ldy
3braiqOSfpfoZeYGkTgISc1Yjosfflkezzp+UBRS9XesMAJk3p3A/HKOnFofhfYBSxYLwyZMhAJ0
C23coFrVXB8qeX8NYecHrOV9TbQ3kstnHBExsNggdaKzMIJv2rt5XJoebQ7sTEuZES2TuelHnp/e
dtBqd6Q4ft1jZ4EBt/oGiP6Pk4I0tPxZFUsR/AkTJlwc+jBkJfvwpHXVTI6YkFj+4b4Vwnw8t9Z/
V7f/603kc/pTfx2PqeRHoAAu2Kks6pzpwSOuKsFqa4cMA4xrAMEIWNW7aEYGiQY4VEu3cwD1GRol
B4o5tbp7aJBL7iLAqO4LclLKpw2fEALpxwmz6RXgSj32nrbEQIEbMXIYt3SHmRTiChzALHic9a8L
KYRvKRk2Ftg+r+4JWaBsyHk+x2C8L94V1wJ833QgeMRkPy1FYMJFTFEFvUhk0VMa5QLvWyBVzRpi
KXIzg8RIfjm7It1jem/ICltUBkJ/Hyp6QKQu29G/qPC5YsXTOOYb/mRc+G/VD6aasxdywbdoYmCc
YMOsvnx4XSkDx3Mj/Gf3tRLKmqCi6/v6Dk7dpRjXKVMKlSg9K96RNwvjLNiYnnQXlKJc0gKMW+z5
qsGMhhZrCUoxtrGhO5Fm0W7rE2UX9Zeans8J4MwDd6Yaj6RSlDp9TTnPIrRyT561/RnxxlQ6cRjc
kB0Io8iu9MW+FJBcjfLRqoyf+Bq8nIRknDy3Q7TAs5OMTFtyuVKdmYJEM2swv0KpGoX+LPr9dPIM
VdiHcYOHoKlST2aM4u1B28BNlVLh9KdIUKK/i5UPMg2kt1h8mQEUyab5OCY4z0VisAIauHs8r+oF
cpXNlSDXb3VIWOP85aX0t/I8vCSumxnACBpPKkjy/bPrcI0aNcxudb24ykee82Hjo5Ud5S6UESiz
WHUQkwGk3wxuXmzNGwYdKoWov33bePdeMIRCnJhxLJYnOOTjhnZFmZGxP6k5QRHl6tHHSicsTEPO
sct9EDBbd48kTjnZEDkJSnNiHhlP8DtYwqPY/HRb7SFI5AcsHzqKnkzN/tJwK81DHep2CPnffanz
pl2eMgqFHxvo7uC9jBGsevtYeA9lYeLWXB2KUVF7DSIud63KnYuBFUz550MalHccWVs68FTlPN9C
HR8pdgvWAfSaZx9Vyi3jck9WVhKUE1pLsDK5h2EZbtwo+wE7dKvBCR1BrsuqiTIdmySS8Vi2HDBN
GX7Ir7HhyxVFem42CwDqzxudB75+6zLhJ1onmMO5LsvaFBVE4knyYJqjT9PUNHM8A+NGUqMNnFGj
pJuhVsYL7lFWMpleVp/qgkYBC+DBcU1JShGYAhzIfdj3kA9L0f7Wu8d6b8vO8KZnJyvmZpMAaFw+
zqWy4nxCq32gKL+p5Je6bPIK/JUVHQMDNJ8MsW3T4erxbx9MaGKXRhz8t7C2rNjkps7tm/KY8NyE
GFX30H85zbithIU+JPZMegmjLySiKlfUtxB1HCpdYdEcfxymm+ypX0m7uzDQ0vCDO+Kf4w4kDQgE
TXmVb868Vb2XgZJv7vqS4s3PCYcbQCVA5MNFZZ3U8DDuiRttim/Nr1pcm1zCSFKWNXS+hEsCMNIU
N0asvmQWtOjFLgWYQIy9ihb893ghpf2//2SSiWY59caXQpJYwtwj31PKmc9dH4+2ENS7AndGcISd
SO8sF7mcfYW1XcwjIcxdbBb0kKhDVYL2btwdRnJqHoA+tT7qDXox0F8YIvfcm+0zkUqk4Go/Xe3b
I8SJcSr8Ffjf+Icpf4TUoMKSw0R48Y5/ARejcSp6qJMYWypQYcdh+FJiss4KDQf1Jf3Gmch3OlyA
4BrfL32r3X+swo0qXTYL3k1J939/cruET3ASF+V9mckqEM745ZDo10g5oegBcFGfuMGE/jECugQX
S72fjuv2YR0qSpbEG9w+U6ZSCpuqPDV0zJokk4XkxKVUiaKcFLcpHcbErHZTEvIfJJIkKbG2+aZs
+O+/ckKTssZPGkdj84xpOKPvvWpMgkTJu4bxrDfoToKYgyXCnodnCBRyYlBpkQe3evuSlwYp6NIk
obT5hJWIYZH/m0eqQ1NbWut37z/ltWkOU7BGjZuAFeb2Zg6CP2EYOER1lgaf5BapnwVLkIK/lZeg
8+GVbD0eND6UPkQdH9IuZ+QryijVtqmdx8EFugibeqPMbApDBJ5s4rmLeMYFWA4IS3MbztyPt8p8
/oWJbv7ODnXIeCrpMVMCnATR1Sx8F2CcdphzZ9TFeP3LNXi2PpLRhWP8eNVK0VoXvFyfmCEbOub4
odEQnTlNXbqyCf1lN/VO6ClL1Cvcw3e41IYzKq4dk/SnkbI+p/B7HXlYlzhpSsUbramzBFmUAJU4
VxPfHWyLsf7UReQp2udBiip69cULpsDeQgdc+09tfojg+Ep5XbbvtEnaQ9t569ixlWFAvPg/Pan3
gezU3bau7A/ocLv+qYVbMcYlob9G5viC8Aw071qatfcEra/gS0F5MRqaNWz71PHA6t7SHrmca5M7
evmZRTqzmzQfjb0tX4TjOdcTxZhjZcEFvkjlRQfztvS+p79FGCkWJ+5DLkF/gHvFNmD/v5VgaFau
DkVHwRlO7V0zVyxV8tqy1Y8PqoGhQQsL/sAZGSJPBPRkt+JDAVc030vvF4CwNlVfxS/BC5eRFs++
XXTiez1R8ZTZsfQ/TJZP4DUOBaQXT1TGMZODWi6td3AuVrrVVKvsHQJtgO9n77fl1LrdQc2b9Oyj
fl0vC8Ot2bV+nVOuTVlsu30Q/9Jw94Sab+IsL657gmWdSrwiqAGcSQpPHtGmpVhsIGa7Ctj27kao
tqkBKEP+yaJEf/BvjDAylu5Y5QNBkLQml/usbWWBG5PmHsowMrTTXxkRfFdIAZZ61XkoMHJ4iyAO
rROGOz6yb39wSpYg6wE6F+ReToMWkft6Y7yE+MyXBnyBSJnU8hGkVw62xSJnAWxkrObJs85XlkR2
MfEMogYOLG6Db5uhwRo1QxMG0oW/KJV8yXHXF6wODfNQDrUuYnTG+WPmb2Qhi+XTG+wCExAnKSEC
PzshcZj9CIKxUt6ftDFMFBDm9w1ka3C7sC1q3wtjYdoC1NHtEverdWXtXxDNaNKzgwynNEx8jYCo
DPG8y5F6wNP3CB7ICIIzBYOUfSGp7vEL8S7558gPWYGHmTjSpBZ0CmBgVrHERUdPWhfQBKVC9/42
04/HbPnluKRGJqeSxb/81JANPmH4JH4Eobwo3hSIpMOy0cerkz2D5fYQWtNiT0BZgbyV4L8nCBvA
QdAyX5grDh986I/YSK86JER1+PPHv2W/DnBnfwxumt0MCYimyS9hp3HvPOwfYO9oEEAmy3MCsLcb
uqTY/F6pdbO4O6JXZjGhLzg28+14o2L1Kz7rbrszg6ZogbmiFuVJPPVjwUcF9l7u/XrOPlLEUwsA
d+lMa7+QFj+qiJNWIoKxlANBduIdnJlW3Ble0Xi1GSla+OdG73Q9Ol2uueIWIcQR32ATRCPoXYdu
2rf7y2y9mi/FG4v5KNzL6yI462ydcK+Y3I8uYO+wSwBIenmA69eaKaGtwwKveKVDrBwKGmhp6jDU
CNaq5QjMu6OY9DWIbFnnnmKnRKYT8Ig97TuzZkhpkL+hthzFNAI5Pf8devt3HD0uyByn2amO5ker
zqwA51PJ6yOufdwOVjJbKSMlW8br7DoKR4N0rrYc7H9LVSefw4Ail45tE4f9w80AAbTPDtYaU3FF
lgGSrtj8gJlVPJN/Shi5wPnOeMbg2v8s9CLp7BumkkMf1ojQei3efWhY65GgoFqG9rjNwVKnLtno
0RGjxzcwgR60TXKtNcbtVcviOKgzB6JAX+J7hBPlVXEDvQJn9cLhDFj+YfKcjuNu/gjhzJBfgEJF
9ln/FKLkHvBwqCUPxfIyfJD8xWkVAK/ahQT/RO6exmePq3zeiQAaDCOP4jssCDcIZ5MLKysWiIk7
cmdnCcTGcjo4NxB3PDNfeXN1F1Vg7zFbBWL06PPur4AiYSD7XF+8XeTj41NnBqM5o6KiKc0UO7P6
jQpR7D562DmUgNM+DXjH1W6a6DV9+Um+ESRvuU9LbS5LVXcASmiXdcwV/X7vs94fSWPh5Qgst7IS
mHFAgEznq4ipTk0ksLs7M/hxmBGGsdrMLFHdbnUq5Yt9n6SgSoQ1JApJ/RHnicXryAU/4NX+ZHLW
b2QQOWYHQ/tF8WBVO7SAbNxyPu/saCVUWNJfNGHsCQFrcOUMZi8qKt3Xo/KZPUKr6pVGlW0WaBpX
UKY5h9LbKNXm3oSOoxmZtjFmhfxUzN+KiGo/oCCZRurRBkku9uGAlSw4uydv6S4/5PaP2c9IXu3q
lKGmiYKhv0PzWnt0Oi/sooLwHpgJa2f+lBHM/ZkjjqXYc5Men0DPnQacB/FtV7ymknMysOIbDjt0
FJiBzc90xagxoOTyxgeudfi9EbLQyUA2zSaV+pfqiUrBdKG2qcZlJ+qtvjCyF2IJtd0w6ngbXPhE
0KrlIgjeNUQAn1tM/zn6hCfxN/LifpjWYz3dmmrNPCZi+zf014ujIfozHWcWjE+kSdj7E/PsMuBz
VX14J48ExlrifezhSF5kHJJzFN34b/Ch102jqboMp/tWxbIK+iS4xaYwto8gVzihl6QfVrRIk7py
qy5HKBGVf70C5eOLgPvf2jLwIxKgvmRec6CBUkmJpTgzlwG1+oWz82l4Vr9KtP6qmOclkAlIXlEr
PLajhzTGlQ9Vzwm6eQXzv+0HNjis6Vv41p7N/pfBLzbQRpkg5OJCmIKgFO5tP0H369INYnOUYyi+
inYz7Z6pIut21gKkbRghiA3smYgSlbrTaHXGZOzaTBR1PSTLnw6QAQQEdM0KM+Ee6VCrQOIuWFE4
HH6APKRbtdJepReP28RIiMJwC2TkSdB2kelqPXWcHuYxpJp0o8g7hFP3h8cTkyN86puDHEPsgdrk
x2eVSqKtmpAvBzyt3HvPFTRmM3VPsGsDjOXeFhRMA2XFw/wqA2yWLmlfR1aILR62ZgnJNBlQ3u38
dIsbj9cFsEKmh89fMYO+liwxJUVvldwmqTbNAJy0tAu6IDMQIK4aoN6SrEsg96HhXOvxkHZUa5Cq
RThtcZWSCLBQemNzmdXGMfVSA5GkfiSsbQb9y3lRue8FMqSQrZxzZmWprBsGwjkfqvSkXGae27Bc
I4Xah3AxaETuaqp3CAkmvejYExyO6l/22tn4qqvzAkABNzskfFtb/cHovPIVY4F7yyI+r6jL8IsO
BhFtBf38+awVm/7UjYEhFABL/7WuPmcd4SjXu63U2eO+fwbFP58AGXNe1un4h8oUqKpyg/fmzoXW
+wb3ibGR8jVGrLdRjrBGFXXx3WFVtMkskjWTxGcGt2AHSdw0XDSz2kAnTb+J3f6t+Ln5wVA5aiqm
v4lQDimRQgepQ/YZZmMTQe1FMnBQrZZwCPZvuLWy8G1jGa6nUJ1mommDbXFwxBwiEbx9Z2Vx3gSR
mq/6GvMNQHYYw9iHMyVMy1R1SS79kIhmJG9apJFxkopNxDXeMkwJ1Y/D1FwOw2F9HuQC1BWm8qaq
mIlouSNQ4WXprGnJrg54bVWAs/5HdIfNUk1uG7NliTQbwgBqTlZ6y1Ogxo4zmmqVjv6uOIkqFNpc
722nssfbnEh4Isb9wqQFh9p03wwVIeLzph3k7Z2tZclx6BPsloAs3HDlC0bVAJnXbAJGVFRkOHfl
x4SyFGchZL6t/pIDnxV5AC5wOABuqV3p+I7ak+GsqaLTn0RdZ3q+75iXxTt7/ZNdQH4qwagBPgR6
mw4RekjyzK00JSakucz78H+FFgfvTvsTCTSzJ7ahq1G74MLWFPlB3kaqa5ZEccQKBuFbE2tCZIGP
yk6P43OqHg5ao5Zn0+PO9NUrqzzONG9JjOXr6Y5G2Eloemr16fvbwGWXaoGgOVKHM71ccXalxE2A
lnufRZ4+9jzYBtHHqxjl+0Kf7d/U+YeZKIeawC8SZn25w8/oA6Sb3igiaNg1VVP+1WhKp1ca9cAH
eUAdxwk9hCnTBEYyBuBJBo1iL0YRJti9RdmU6SiCXsa1qvSCSdPph64m0zEOnyzyO4OhDgCGN3ep
JKEBFE6oggMG3M9ItC7T4Xy1xWkKngUAbDFdDpKe8nd/kxIpfzxcJQQDrsiP2/kZaU+/wRO0jKu3
1bBh2aggHF5LJ8zmJ1x+oStTWcyri2C+U6qoC+znFI6VhN8N8xcHwiMkMoqFaC8FDsin8567Wzgq
83UpV8QHrEWS/qFryU/SG06ioNwmJjR8Nf3zyVCmAMqshX1M5qgnxCLLGfQE+OcMI6CtTYCbsVBR
awhqUTu9JJbHZA15jxuMLI4wPiXmOfzr3OvJjfg6zyUWtS8p6u96lIb5mMsLCaO/IR+qMfCFU4pd
QTjG86v/bX+SpYczppi3eOgSGrZx+x7QEga9cC9EJrRXsTiuWJFMFnYpzM0/nHzLDCRgpy09b8Oy
FYTqHckIQ/r0dyGkmrSjFNxI/hf5ZPmzfvKZJcgNKtI/PPlp0EEW8cx3SBQgHeppu5pJxuBL3tKp
od0/aqPZnlhcsFpN+Kf3Qr/pzqdjWhFClgY696N5QOetCRvP5OAfwqkKl+s6lDltVlIOawH7uyXN
hqYs8qmnTruYkXzv8RXfDXLFWuLo6GpoHHvAQjfZdYczw8yxc1fxolqWgfSIfNSvxJVAMBXIbUn2
RuWlmYdnoOu+wiCTEzzCJXWAPkGiQSypMcWJcvyRPrLvz6oytDIA+YRbM60/ERvhkbIrg5NEbdKm
BXQGwnhK9qx0qaCVGCF+skqq1oSr1D/iYowyBW+GILhr/pG1MMZyt5NZvpG8Z0lr30Wc7bbqHmN0
Vq9ba0hdYnh7if/ghMFfe5aIwYEktPBkB2WzV6z+mkW8wI2JCcIhOlYo0D7XQ+7YZxAXSvy6Q0do
1U1Pp20ZS4fKjPDBS3XVoAGxaWFnRQE2yOaEZtGS/kKdH81hxLGOwL+glejuSUj1Q82Buck7z1+l
Vvwfun1zeFKxU08OMW2encX2WEakSdNqBU8Ol2jkot8yTf+XhdQ9stylU4rQTkM8/JVHnOKwyZkb
wkcZ6GYfVtrI5R48S+cTJ9WDBMuZdWDScFX9picjAHkb9IU6ZHQZ9yv3vvkckvJajUNH+NxSCBoD
WA8ZXzYrAyNkBl4nwloC98cUS1T/VfZH+8yFe4hW/r/onJMMEtfsUIiHTvhAEssau+/NQdoI43Qa
HuTixZMW8irFVODFT0WINyhK3rRdazi8ac9qwb2c9z+byuvtomk0WnzlwnFbGn566Bh+SOXRa8KJ
Ad+88ih9T7iA/GTRjZeAbkQ7PgCGrn8OUj91PXS/B0Sntjcb1604Ad/4HR1olY46vrIWai0Nujdq
bc/8XfG4su3Bt+ix0a2ZVW3ptdfdLcRcO57sFhKBD3WgqS2sgnTImQ3exgI+pfYC1XytlqdRxcbk
bn51iLO5sKigvCyj5eDdstuQCkXR6IrQbobqv8SUZ09yezu5k2FtgbgZ2c1n/SFv6X5SGgqsR4G8
ANM+P4LSdubZ9t286w7HiJimbmbC6i4lNNib8hkI38JPgJC4/TQnEjIP907i6hxgP5jfyUJXTDhn
rT4Gr2EzSbwRGk4P2T4D5Ptd0V71EwKe1ywWnQLTNcppbFH3W+KZnZFJBRorzcMwjWVpfpGEzNAT
LHEdHc9Bjas/9jszlE8OYh9Qnd5jS7LCWm54yVREH/gbnHDFNivT0W6KbPmuo0P0yUTht5ucBGj7
6FnJtq1PpVOLxCjeCjE3Cho1/G/U9OddoPbB6/bI/molZ52I6gFw9/TylDW6z2nBfOLwmGQoNkFS
M/ecZW2jQhMJKBw2Lm/Gq2XK1i47A7l6VWfp8wU+9rH91Mzf/0hwAe0iLjEMNb/PsvK0X0f/gHCb
LoX9II9VW/YOzfUMSqKVjMtkD6umi1FuyNfnoLV+46nikrqNjp0RPnHsXiFeHOCFXOrq9sZVAq83
R66TzoRYuGfDy89Ujnei6/RF+AiTYH8womEKyr0Y62wxdbO/dfP9/aHJe5Bw5fYXKahklY9Z/R0V
IdGIPGxlVWbeKg9Y1olGOMcY2j6nYfpORN7FXhHb2M1KaSaL/jMfmHIvlH7j/o6kHXPOUnTXPYMN
LNu+pB0bJ3nlCikOAESEDZBoVpwf4pV68xeZY4QR3FALBsfTOqJL7O+RzqB314W5IzSTOTmRVhiC
Dcisf8qbMA+oKZo/Xj9c6m/WalABQ4AzWkdTQeprPzbHnrt/dNZ/JkCbaTyl6QvRweW9+/F1jBZW
m9vCY/8I6kPjI1DINLTJwGDtSTdxgekGERmQ2UvyeXBHeQmkGcG/QfpYc95mprwAA+pmuw1/8P3w
TUqHhyV2m2Vc+oSXCrMlA5AqmmzJ7MQfpyfkUSQv9aqJ61zCrc85LkLF370RweZFSCCC5S4R2/XI
7gEocE4wVTEEP8ZAwLZfd+/AiSmSTCEvWP/AkVAIzfiQHUQCD0EAWeMRoGtuOjzKnnNSgk0nuLiy
eRqKAXENCC/WGs9ApFEBTXZjLG5/dtdIv+PHOsyuDu5nv1DmaZc5PV4vjAoeNjrilOwKqHaT2/sO
vmDXCkBctg/QpQSzSMnL6lvnzjPLqMiGoDfrLwb9+A12ASWL58Fy8OgYStx54n+9oc039J2JxjzZ
lb6H0pbzdj2ZatAU12HvOImel8O4zA6DQ67uJHWrSmVfoF1SMzlOfgFTv+9eDkKGNSKABgPzPRTh
U2Z2JKpHutVKrXUtg+mBjmeZvCIxlTIDBcBldxAWrmVK4ov7tKOHMTGBhbfuQEYnhQSPdOf+YNf4
N4yOp7ZYAO1e+Li8kvqaD1feHcF8bKH0HzEIZrmdHvxQbmvpBaQmkEhVwnhcqPKmL1w0wF9EBdUG
Zs3Mi5Gjx2A6bG6qda51oXHAzbFrxOS1jS7tRrBDrHsBfPhgWOE66R08OXcda0bcQGjOa6lcqsyY
cBGw5a2/SrulQ5RKEALxKmOUIClfpEmOJIH32m1zZyuvkaIiIw6v241O4covZX2NpYOGLrysHJAj
wNKZQrIk2QHViBnIE4XBcopDHaSMZKgVkTw7tNTu7aHgt84wuFk3TZwGhVHMgCvLQq4EiEW3GsRA
kdRieRR12Od454ML7EwBko9LFrONRz/v4Q+N0l95iL6lD8ZhYY3ICNnN/2Wx7EBhOCS/OkhjYo/e
QMID3o2eAFV5Xi8h8B9ENm3HgxQNHLZIb/NptWKGnmZocMbNdzJXNzqyMmmAhSoTtLe2ODdgYDBV
hzdeH00uS1Rzo3TYvh8pkwsrQHRof7tA3CRD+98d2cGXNAoxOORX24+RpRTp2sH0VIUoQTvlQaMu
yY4Wb+J5JjG2SHhFN3DD/VRctY6TjTTZM+/I7n8lkGGa49t94iUoGQohMInT/0Lhc+LuHrda1IPo
D3+FBj9uFWr9hGrbccw+rvObIP9CuxoASEHwFOVS4TAeriDR0zSzMaN4wcTRpAzYbDm0xs3RlhT1
e2HK/TztEoBs4cpaIot3x61sv7GWAkdfkRRcLYUPOk6BZ18BGJhcs0kGvL6hL0rI/JkuwoLyVdxi
DB7jpericgtAVzD4RIsCSj7hMnj6vyUQB3XUTsVPFs6rB89UVsFCKa1Yl7hEqkkq8pMqIT+mghDw
XKi6O7GoKgCouDo74Yrlzkw7X+HqtdbxwMhkdTEJtdquwfHB7WZZYk2Tjc2LcBkUIPDrw7xFSk+C
LXao9SS8GsNS4pY2LtJSP/ckbWxS1vHpIF6jftuPb3skMgjA0pofJq/NTdfz6h18LgbNOYqzRyx4
gKyWT1DRwwleg7pYe25x9LhQsJU+RmtFet2gnpKmnrvA+6/Y0PUpd/jfFn1jRhI8v4b3Fl+au1rx
BZFVify/OpvIJqldwlr6cZk4RzJihjeeomln78gK2nvkPJcUoi6kZWbPRRiF61TSgrBO9G+kvvCn
Gh+fh10tnd1UmCjDhsjiiD8f0sfVu4f5Xbp9/em0WBucfXo1+4phlQxY4SuGpfegmMiVZ75cx5Mb
AH6ilRGaJsdnd28dwvw+6pzHl5tlzg+mrHq53lAU2kFCXpDiMnk6grmDwICvx2yaGRneLseK/JyU
ztxVsVwvaV7hVZflGFtN+LaJSWe3kXrwvAVBg8oNVCb0BolhJZgtNtxDdALgEstE+FI9eoppGE6l
fwI9J0OES2IRbF3A/Atk4GgcwlkBJ3PM1SpPKIONav2EmVvwrXWtPtCUVAItp0eFRr0bRpgsfAmx
8dfUuCn+hc9z2uqC2pM4pSJiM0q4NL3/eyyC18Il1/Bn/Lo3FHEE5ktWYodWzL6Evjrrv6hSIbJT
3h+ewe2Ocw8h2Xz4TzIpxCb0F3SrAxPijw2ywSorUE/eBpqxRt1oRCL8rYMKCf//zF+nM8/tNqLw
HbJ7/zbGFffss95BuAY2b1Cz7CcjhH1Fqv6emyoo3OOBc9DHHtD5OKJxmjmGekFFWNy7oAORh/yS
Yopu0mIHr7PYw9cD/HW78wXL3YAaf56GNdC1UKQg/uPo0YeUsHU+mjda3XH+BZWvNE6LPI2qqm9c
mYdB2FsOdOi75rKHpRTKwYiRwox+bNUiQqf9WHx9rVpieHMYWOz5XaVm359tFBysoOwMcu4JAxln
lSZM/h4DTtAms5Brma/58JrGCxfQyQTx9qfrzTi9/Ik1Yuk5SzPkHT/FG1oWlEsDB2cw+mmXo7bd
GdwQ7bPojN+RVRWN2KobhXKXz8X7BMsvOSWeuH51R5GPXenQQlxsr7cW2/grnaKO/h4qAWvHzyqg
d7mitydG9nAjP5k86KWXzYPG8XO5pvsvB2t2OiGOv6PqYo3Pokel6LsAo3p5L1oFUs75TX8y6dxC
nscIMpyyZ+zuB7VC8TlcjPI8XkB1G/1qO0OuHPvEFo203vhRUa+3G2ZT9rRMAxTGjnRgxJwlRfAm
13qeUPnrbVVw5/U/u2ux6j9sPK8R9Hy+enC72pr3qxiiQuXW+kpzs0qPnH490cxDuUA07vghpNQj
eHI21KqpEn+jZn039WskEImS/TVgVbsvht8zcmaovGGZ/GCmAc1yfRjT9QYhlxot6jW9cKhFGXlj
53RPjzi4EmoCErz5qnO22fgVAobuY8SDTNkleff5r8ngEaiJREtzmOeeF4LeeoJ40BvdOuxM+DOA
aXNaXLhX7YzW7smq48EzDMBmTiJnvnkf8D2l+AkQ9Z4nbzLV9AIISEAHdXN0m9nhMHfxYjsfXdFM
HwEPGIvA6pzAvEEtcErqdE9WcfeaWn0qmEg0m9vKtl6/eY/M/w5U7v0sDxVgHnyWZZTDOUfiQpYq
/UhEYO7FINMzBUphuS5ZARMdhmPjsav2KhO+IK4GCJuYmIKGCZ9ewqkWzNJ5+3fvGhqHpaC39Djc
hbD9dKsMb7MIixZ3j7EO13pz8a2xME1FBgZz9Ng6rHiuzujIwZmRMkXplScuJ0kxKOGCqlwq9Lbw
PJzXKfctmjoDxsLqcUmKGjzwJCDnBc7L8Ni13ZWkoqimxK7CKOxzcvAFzIrl2cD1TjwqaBC3xlqm
fvpk5vm0mRKWlg/p/ZnIgp9JrLQkJ7cvjuyohL7UFbfL8BQVXBpEC6DpHvSG+7sqs5S05QTwVfYG
QMNVchglk/kV58ezGG2ICKDwEVDcqYBKtTyHSA6oLZS7joWWI9iDmOo175v4QJ+FAMJYU6SeYqld
LqxfAUsSGTw4uwmmgKb59z10qZoGUq9IMy6o2l62Edj4OAoI2DBZW5RXGgZqsZjndTnOQRv22OBf
b485xjrbSgH5T9HBSIVsKI2/1vbes3dSaJPxcGwS6hciFpf9f638Uj5jacy99BKbfgrLl1CmQDLw
ePunZ+biyRPCNqMVuJO06oPOxZozEDM2oelfBCpUiQAU76+7ozZF28XAzjWh8vCTTiVW60NLBJwi
c6Q+mkrUUH2N4v7fINcc2eSXV/80jqyrO3mKcrW7jlZc5o670lgkq58nXUONtWZHZX+fqylEsMuT
iG4rrYMzTW6ajHTSexW292MQUCNjkhudFCBA7MTZDwkyjXAjmB5teAqaffFFBdSym8zdFHxFQzUg
GtVGu7kgYZ17sySna6Wr0gMYXPqVISS23YH7A8pMpxBUaVuJBMlmBFAn/bQ+oGB0eHAToUhx2tMh
1J2PW7fGmyzzz5RyClYw2jNWVaV7vfjRlrE+eip4A9wbBwgUg2rOVWTzEDk/5PUS6myzoV4c6ukk
8ISL/pw7eV94jThWIQsr4UP6IkYbqN6dNp+34+mjRPiPdPILfdDcTjAoNUg0wDgrywRcTTECUUT1
zfFALYkGf+5QDX8eEkCOaNnhq/R7WlORqyYB5kPWD8CsyI7/eAYFbw0MHAIZb21g5ybrAZyCIc3/
HiMWTu5Hbjs4RcBM1fPq2B9jYSxTlRePNnhmAHDK84EaZveFt8AjJwunvnToViKR8Gggt1+yaH28
IRD7ZJoi91+BeTJ+Ha0zmU3nNUZao5O+Fhmx2LJkt/nurtcSkuM8mP04fpc3boQgL3XY0XTTc77a
yJykOUHjJP644akNv3WAziBr+hBOsPTE0E4Npwa0FYPIdhNFz7jRcM5xyzxIMIUb6+x17SseoenS
JaAMVyxTAZ/Upy2O5DJwvyHjkk6D7bpEajC1wndREWoL3oK5DE++jMpkYgwDXgMbyqJtEZJQXfLa
Uu5Q++eOvyN/Qqqw/N2xLXhF+bWxBHETwYwagagaCpX9CxMHsOOCOUJpU5zLyhG7Oqryee9n3VJP
JS+83Uj4q4r07DWku+ULWzelJyrvR8TqOoj54Hmf+sYTEhQFle3EyGTAZdtgUT4FBdiW4Z8j0GeC
odR0L8n4VYCQy1ytUEb4tAeQm+JMViKjwAbW1br723Q5viV2Zy1XNsrf9GvRAQTFpmvFkTpg7FIu
a0wVCgBl8gy8n+oG2g5oH2UZ9U9vLepsAKrAkaN1sUQY87EWO43TmIED+4xAxYiiBlWLCC3orxDM
MI1IMjZcX92Ltpgi2KuT5TXuDQAgT+0VQ8suUGbq3Aum1z1XIlexbYcGSXawO9mEpD7B2I3Kh5pm
xFxSPwRrcZ5C3yx7GiUrPrUwf7/DWNKvLZHhI3a2zKEVzyOdY9LALrGsugurtyIBbrE3C15hyZsI
ZYrGR2oGkVnsmGnQ8yJ5k8qewWoMslZCDODNy/KlZrphthxNjPtKOvURNhxprMs52PZDbLMM8PeC
Uc4zhFWVQk6oP0S1bUzOuCkc6kN8uE4a9QNrxQKEwCUIagR3+wWYTFKRyd4E6wG+4GK7nYctMDFJ
MhbFkiIlmzHT5RtoOuecIczAqI+UwyqjAYnncO+YPo+zCskK4d4N+PPueTCBDSw+Jue/+ITLHL7Y
UmWkXq2zxHy7dS12WQq0QzIRENEhhr2E/L4HT9KmjEj/6IOmymsb2KheXySvgWPkEvfIKhAtGI/u
JZcWX2HWWCnJ5vEhq1ZjzxgfHD2Z9vb46+yeUlLYDlZ/YQNy4xcDlyCUS6pLO7A2aFj53JQlR8j1
mdXnBFzGNyDm61kFR0f53lQbofDMcssqQcCMY44AE+K8450UHzjzRkn3Fzy9qQMsjA30Lgey1Kod
7AHEgBMXCoxzuwL6z5ToWpOn1/Bh+pxBhOXIvJOuRgYn6+Rm2E4/Pxb586aW9PeelLSnt9xEuAFj
LmtjidKec0xg5AgCEtUQEG8LBVwQrSKmnHORKfMKLv0L1ZIDWGtRIihcSyRdEAPIPSe/nF7P6Izo
hthHNh55GZ87bmW28F0hI0Eft3uVSSK1gIF3L/M9WZe4Wm4OydSAZGIGPu93i1C1OG6nrhg4jI35
aLtGwTJyCG0LDXcur0ToAjXH23ivayfOc0Wp2b7B78DB4sjF71YtfZ61JhA9D3iOfC8DtEHutpVA
JnQfLzaXAarSU4J10lW14vcvnxhVdxy+/fohjCyj3pobzKtlmPdY5+z6z1n/p1XrDMDqbW2YHzDj
8nZvn4vZZf96LmfYA3McR3qGL/ddN7NMKciYP22iOmylhvyd3CcUsjrCD+rg0CECHglY7igRsq4T
WRgvQ5PcR/QULcXdw7Z8RELzslcQMaUQZ0PQzo61V+dkRvvRKAxP901LWf+2HMT1YAiviMHUVymJ
KbKgUyYDr48+Huf+lJewZpyZw9F8Z3RLzOobdmqF8E/Yko3P0zzU3WOYi4VEymLXcdQB/QyLG2YP
e0HDx2hQTccovVNXzYamEJ24ep2FY5fmOBxw+dYG9Dh1t/AnfYL8NKb1ia7tzz5O1gH5zKTJzvdo
8JU4uyBE3+uy5zNs+WXHYIgvza3KYu9oejLhPYzaTPMWPX0siM2eOR0V7C7HWVq/uX/0rt0P3Z/V
qvXoOnWmS6Yhy4KdgokkJbbf1sYeo8cthhTIIO8Sn8P2QJ/UX1CWnNTO12iUf+ihGVm5pQTQ5xJJ
2LP8YJAp0r905L4DjrLFKLq5w1VXfQzYFLpoIkEusBr8bTHujj9v0wmIg04A2lpUQKuWJlv1cQ7H
DoPGNrq8eqt/zH7vr0H7TDc93qFKmXRUte3UuL26zZSmwcUbWIxdCoIaslZS6F8z5dCWBPB1biPI
34iN15KVyNsKZKL5t4M3mt/YuTBAj2OkRDlHaPChXHndY6eMPRxiUL8nTCRCfAKGXUqMZlwZYhpg
7gSCmBJ+7a/6a3/wByFo+qTXx3KWioic+4zN52nesmhaKe5/Pwjdbhyzq2vni0wwpcHPJsgCgUp4
pK8644YEyCXOMlHeqlGV2cNEzBrxg5OZt8Pm4b7vJw7H9aAxLDcOwLiIb2TTaLODDjlk+/miKjdd
gWA0r7hT0WmBw10xECcLVE8Vafd/6keqlzRS58jv3r6jA2p3eG2c+giyyLBMZgF+LPcNW7eDw222
Vv1ene6DButEaMy4Dr+lOHOMPquWG0yJiajkFUBMG7AaM1gbslFmwAt7xeszVFGLQxO1YE0StkwH
zuypAd4oiyE2wL6tZpxO0IXpEharZ8h9K/OVZdFzZ84RtY/nznqBGjBtiegI7zSiaMqz3jps/oEU
eefh7aaDQD+fAHCkoe62tvaT4GJaRAF//8BpBgq9nAIQWTmaPA7zdgMug0Zgz5PRVyfGO/blOocQ
opVqbMq/JGhJe1RMloRCWx/kxGTI2C8XnzOP0bq4MivVchML77CbSRhab9yRTPWqFKUUh8iP99pJ
m9y36hrqKbArXDNVNQHKXTe1B1oar7XidVX3LYqt9pnRMxPHCjzjL9ja3TfLj4ODU/3pXC1/ZeFv
bHQuOSLr8vbGydM4VZehFgRSliqh5hr/0d9+CLBP9Jmi5/kaboX4e3Ck2uqTWuv46M4oAiBzwwXT
patgQJGrN44pAt9cMGXp1lEWq55wrc8Uga6hKH/NRatVr5yJ4DmsI9IIf5Zv6RTV4qXGylRJzSAb
QliphS8yFGQxYAPXFNlL0vr8Rebvq11Dlg2gAfiSKJtRZrfZw5MThb9QasL1GlIwv342VswZ/xKf
oXASXO8cDKYQRRf7y3Xp3JVG3Hl7DMiBZhZ0lu0pRfQ/ij4uuaTZ8o2QNBI1fRA9QU0SrFtpkoKj
QizW+j1QjcEAO+lBvZZDUvbXAuw9nO99rLRj35598HAbPrTovDeuElqmCuiGMod0JZ9zzlTa7yi5
K7c2IOJK4LBqdFpBf2mDOTDgQtQmAYS6mlCsF7GkuCvKB0riTiG7IlZ4/D/dd8iPPB5av3wSOfKb
anOPx9sFpgZ6AIuv+6onHQ+rbZpEHsDMaY3KIPoJGo9XFF/RNb8ShDDMTEo5NzqGe44YK227r61S
XMAZIq5lspLyYdxGA5QuXvPcsFu7Acf/D+TZsfJ52du0UAlf0qPw8lHV47ACujRY8lsg9JiEpjq4
pr4s87eGc/izgGqf/Vo9FvANIMmjHy2KqEOWxSIOWbp7Zle/I4CZQR74T2u+WRrgqNVdhsLlKH6m
WtUSOU5pl2IEPJHpwGW5JuRv/1+xo11YLqLzdf8xpYYBNWr/TiBskrNgCy1U8g+uVB8FAzXqGD0W
cDj9HH3p2kpx5UW4VkuHQSMhE54a4PhziLTg901abWyntvfZKaSgBVF+/3Tb6LesCmnRBhF9NuEL
vhi9apQdGoo7zpkn9MkkIlUACkgADuaIle1F3qLR9tgmn2Hefm8H0JH96uPODYBNtUVWCP1l3bQa
8H2JCB/PJqV6kJ0ejIYk5xbFY5Qi0+EpTm6BixSCioAYExP4zlF1uplytq/lbin8Eux2xYd0PKV4
99CXuB4ZuwVexA0ziLPADRcopXiMdg79zAAJ9wDDmSpFTtbtBk76Eq5wvMya80ZFUSXEEceyxnnS
0ueoP6ytcd4HlFeak18ThhhCJemWOscjn63o1IUdYP/+2T7vO223k8sJ5qZFQvTJd3RdHqsxCT9H
/hsAl6VRqA/APjLodupweP6z/0LUm7SNp9FE+gVdDi6//rf1V/J5ynTSTfrNaJnQSVEr6wF1mL64
JWclqxbrFUgioHYuxEBOc9UcdmI6v5N67eE9N4TJ9khAn3jCZSxXOIIFV80vejCU8EEm9ctGDNQG
lbqA/5T5+O8VbZ5TuyNkhDV0Kg2aOHHVP3tdMDDqF9DtouwxNOlBnPDNCzqdHVEwbXOjwOQE+gkH
54WRyhBjukP356StR3HlcsjOr7Y1bnmG0EDb77awYoFR09p5fQxtiX/IhvnBkNGxAbaObH8uIEEV
pzTsP/fUxvl5qlQkGwTsQvFYf6bxouKGVVhVB5W/QtROGS3WWfntMJkkQayE5Maah44tfJLs+NoA
t8RoNUaQxWs4+DZy6XtcZwRZsFjrrhJT7m/78XenprOBCPJnofEdX/lnMGzEIF3IJg4hWj3mCXs9
SvJT492JRQ49Zv83+pzpiAaUYzxLhuM+UvRDX1ip3kRtd6BFZObqXpO6K/94DtCb4JWHh4o7Ck/D
673GPhFql64UxrnGXiDCk6HmunfeKSha9+Pfht0w6HO/ywQWewVxR4tNfpTcrcjps3Bam2tSnvsz
CTLUnEyp00g1l1Jk0+dx94t9sZef+5x9WQLCktiwox76L7Zi7E+4MBZo4AQTkyCUrLTsbs6oOD+L
T3kgJ1MJetAwA47NDIw961+DIyVYyvkgY3Vlndtu4sFnpFcceNmxjhW/RTfpP2xIxLlRRR8JtK1c
wb8eoji2e/Ep6PF+bFX9QJBiCiBdM1sJM0lGRKBWw802eejGgH6Ehm3sRZ0amwhCEFb9M2NSDJxX
o3EyPmJzn2xHXbIq91NsIu08VKlzi+/LhBuKSRFVHZgC2qIQmmL8SjpGimMoIoQzBSZVMZWjKHJ2
Thk/yiI7Cy3Pnph+Rnkv03iOn2u0TRjShDM43Fxgt/XLhivo+nMLEazYbSZoamo2wfI4VI9A4dkt
piP/NSaoYExJ3Eisqiu+MhVJ+sftfvGOIv2o1kMTfsnORtlU7VaVLbWkEmAxeoct/U7zYwSy4RPP
BwFkrea1urny11t9Wztnc7J50NfZ2BCcyCKFuE6o1gjS1IY6TiPlXgjsMrWdwSiHQnjIkFgkrZ9Z
AiqbGG6TS1MNnVzf8MSzlmmeggmgqBMTBnZ0G5dzV1xk1u2xzwnjsrA3veZ32RRuE8A6js/VSXXF
UzyG5C8Ce4twBENhd94P9HwrhaIhlqx6J4qpBGNqmTmQWXc9G99UIMjxGZjGSGPGbgEg36saNRbm
pzCTkmniOzrchUjQIvhM3/tBaCJ1C1QZZg5IK2BsTvAxClgC9TgK7Y9RJLcpBPQSCTanwnBdZ7SC
UogRypXnsEL6ur72f4J1y8MAaUKjcJcdrK2AQbEc0gbDA3HcgcGVBgBHGZYE1Zepo+CBRZ4DQawO
Ip3kyOGhuYUOJJIvI+xmuIfaqv7zZwB94Z7pmIGgfV/P3O9JLIgjPRVzz6GUzSMxSf+t6MNY561s
y2cyPgH0tndts/wRkGBfJnupMHbO9RgTC8lokGVw6aRRPtWaoHSxyTU+WDUhfXSRanFQ9oT9jyZR
MUYUnbuXuBmTUXfbMekDw2cXq3FOqhyLM8vKRdTZscMPWPfR3pm19frnzdUXhgr0qWp6pYCnWOrc
w+jjCQ5uKbQ2UfyqNGou2pkGsbBXMMHCJMWpPDUb03FDlFJSefVMxbTOcY0wmQT5SrHes9jl9Moj
JT+W3c/FHX5VTkh7MyQJ5KyJC97f+6lU2tTVydBoDd3EfSZarzvIIPYtVQC+Mz3G6g0Wsd2kyOuV
FBYoulx7touBk7Ilka1Fw5vRTRyI+Vi0Y7ZieCSKI8gTpr3HjIHfpPTABWY1p20NHAspexJQQUbY
B8GdO6zdhj9BAVaCXkPtC6gOgM+rZb/CgncvzmphN5fGrqkN+5uSluA/o9VcM80QQgD7USqCOBnH
J8N+TfDKIQNJWATljxDLGC2DuaBw/ilwlutBg+B220lditzRZyYl0EOp4ZJvORgW/WQX6RfoQXId
XgKO5FTYSSHRrInxFAX1nKwCMKu4RHBs2ZI1S1RrQOHagog6PofPVdLFt0ueSPd0K6suFJNfsKK0
Z/Bpi0sKACZtjtwx1O4qSvD5fMhcBecExKe5YoRTkeBBSKKzJEeyeok5uOO87OEEeTJeD5qpfriW
PT/0gta4Bmv4OvB5UR2DHtB2DicPr0mppv5bQDFwH4TqRmdyJICU1O7cinF3gJYloxg1g8/lB5cp
B2tzDJyiQfLq+4MVk2iqIWMQlFILa7jgRitp3lQf+tiICkw4G2wv4WWx89abJd3E2WdLmKfK+wYY
UfJnwOaPN3BLpS9ew2CTsiMIboe6rrgEXXFuw/DVOd4L33GN5/z+So39CR8FN++oe+nMhsqKaIjz
/SiUvB7RLYIGwFW9rk7uu36LyiTzW2rNa/A4YYZxfz6sox3KTqTtne/gPPXqA1slRaZlUPVzfUNd
6VEJteJTvYuBsaADyjm6DWjFfZEbUjtQ+wdvWISzWD/gzSc0AS6vLASzss80rs97dTXlUNPMrX88
/y1SVZ0iXTLX24y+GzUrqnHioEH1g8TlEVWluJBD9CqHGWk5YnYrzaYRuSnBL+b4t1AD+oTDLmPM
Mwu1F+S70BI7IFe1xjwkO4iNfXCAPna3hbZrh+uXC3Gtj6at4pDz7RauqoINMrivMhKvih1csJV4
MvGMNNoEnjx4TcUJ64QdcZRyIowQe6nNnYOdedJsT6P5jDe5+2ZklrsTUGzrKoN+8QRQZ07aEQkX
x9UZV+fNIkcVcUmg9TYeHD5I/w4gP5M+DwDSbbpjdFdc5+r875DImXLpywWGf8GCr8QbGlhP59a5
yAG9k7i6mfScKMyM3Tahdn27yUaSsHbkTdL3TO/K4VPMci6CFL1faKiv4wWHbtBYoNlDFAmyxU2r
v4IE/ENMFmzC/dD54Dp7JM0glZ9RKqmRBt0AGxuKx7cf/47noB+kuXu6rWLCYNbeAMsxNHn1fkcU
+x+Vvevax9y7olmimzGzmxZP3fpcCy0cBMRXNz/J1Xjd0yBr/ZsFw65HQlW6HE7O8QW9d+35US1A
DTVzEX6JR9mCiXcwhQFZjiFyZP6xNsFJ61ohZkz7pYX6XxkD//8mvZQq0JvbnJbrz0gqm0l74ecu
5HtiTMO4QGO6Mk9g2LLSKLPHoQY4sttby3oo7zloTqzmRNwbLK99kLOIQ7aemD53kJvYBjNUKELu
+bWm2GN4gzj1w9qt1d+cg/JJG5PM21czZmEwnLBA5rDZLDPxWWyV6xnLqd0B759s1FO8AcgkdcBT
zZeg8RPr+Kz+EDqsN/Ac8i6cvbLODorGEqyfFK1qggteMeMQq3C1H1GXSUpe+9aNg5jvTnVzckvS
utxfDVKj+msVhDXKf7QePcV0zK/HX/TQ2fXATyQ1OLKx7Y8nfo2VgHnabddICRZXx2Sw7WVX4fSF
daSpke0ONRomsazbq8X1yNtHiQQp+OqL+7erDFUU1DeC/xyGi7UEcnivkzQEwovDzLlS82VWOdDz
rByV2ZLSkihQ1Ed2x7CkjAHTQdLAmDZ54Eq2r2ba5w1pQzSUGnSm+76zMK6ZYdei8Z0tS/7wN8i1
pq2CANDPM+o3jS5C/iK0gDT0077y5AjDkEeN2+LS8d0Q94/1kOUyd0P4bnZHsPYAj5M9jiTBmPlv
B3eMcaVYnRaKWqP+2+09DDlmU+VmzlomeW63ysPQ1AkbNfr0rEEhyJhgHoMo/0stNDW3IBZuexV+
aUO8FMFhsGXXS/h3oUXUEJs5zE9uesXV4OOquRzBYbflacfZlDouxEZGvssQIibzt132JA3qVBOm
TAaA6/Uz7v9BSVgSsnRd/JH7nVJmrP7sJuoaHfOY/QVZ5V04dv+d0w5DG/ACXx6t8FFJAU+s/cBl
ZD/H9sFAYlQZbd7M7vYV8HmyIM1LrMK9UvkANavC6mYkYCIu3uPath6TJgEUg4QxPTn8QqWHK/Ro
QArgw954o/Vm0IFHK9N/RRUsxDKvfddUyHDdZusDtH5Q6WXUWt+k1hXDSZTbtJ3ysUttl8ZgXL9h
ALehc6J6gdxk9vXq1Zz521Yt3K3RAKfEeMXdr1412Pway7IaNRMCO64QpUEVWUaKusifrKuVKjY8
FYWOP1wmJLw8ptoU/B+I5XBpKgi7YRjG70BGZOSiK0dFPhT32VfFhk+T9JkSiDLz8icwOcanmmUU
QvKPuyE7GU/dQD+faVqwGR+JLTXE7F8O6cYiD7JWWdrcqehd8V513VVLSx1mZdWHSP3ZVGV2J7xK
VMqGxJHkenNJWp1pa/YjICHuWjwrqMc0frwYDQbEbX/tcmHh4dxRAG9QF0Vdc7iGkevFubAwyBe5
keSEZjHoZ4gsFtNpkqZ4Lqg/3NckUQJspypRtljfNJPo7EMJ21iTozO/H4buliz6ED+sxYxh0bYA
H2ZXHld8O8aWH1Rxl1cWtdZXXt/9UrgYdkGd7fngtjE6eSbrHR527YFmqkrUHKWSG3p/4wTNFBzz
Pm4WE7fnojkC2J9vTMfsZlW1udD/aeG8h6oG1dMCNiEkeqIqRb1cC6M5OX3nO4AEG7w8RkwVOhq+
OnvV+9FvDSEWBo/w8QVrbDvWXZo5ZIwyCZb5Axg8/IJb3ZecZWKMqoIJfwl4sbpLYpAeohfWkkA0
l2G8/CXWRJSRTFYRfUsFGXDXg90M/eOn5+OEcXFGOzBcWJ4VUn68xBEm+xB6zoPDcwABsGg4fOUG
IPYyA4YHzxRXpSS0n7hDPDtOIVCYRHQij9/XWbQ0PpiJxUPouTlk2XmNfjdRxMEgdLKyW3njCuws
zzWK4Ti8kMajEfHFoZxJa9YxtyRtr6drD5+6Kq4M0o8Wx7twRcKN+5Q6LwyJVYzS4KnXCWtw/GuN
fD+SDGzQsHk5nB1nhrqTUGmm7l00r9TYof0sn0OHt+bzJpDxzHWKCWxbuiimhGKVaj0aZCnjcEmu
mMN6DQJf2Sqb9BC514iaPX7IzdrMr+xCUr1gjW18lcobcz7VmLUrbmm2XDynxSS8IQR2IXH+x4Hp
6LjGnpNpWGsZl9zr6zDaeZGJ8xqSanhvu2lKi8kHsylWKa8Ep/qbxzz8JgZWOLdGOyZF42dyX8Bg
xKmfYQKmcRlG9Vcs56WLxV95q6mQ5kYvRQt35mBH5CReco1PtQ9D+cxeLC3n3VicNzrBp0hjNrZJ
KwzYyswYNBnl62INr/8Vn7Kv9Shdk5+X8W4siYLHaVTQK5oh+fdusdEW5b1XZIqt8D77URI75c9q
xGW7r/VOEtkOhHiU5cCx/ZlVzqz+jMxdHzLDTqAQ+6hE5G+FAOMC5HucTVATtjdY76ob0q3hzPPv
qAAvfjBp8M+t3A+VxhES/QAnQoX5ISddjdeKUtTLPoYXsOU1CyPLrFfbABe/afsUCbEJTFZPWUdO
MNdMHD83mtbQ5z3/LRJFi4nXsAryC8m5Tne/4XuQMuiaHAU842lo9v5a7mblnQVxhZsUGrGRuarE
YodX0CqKSgceDs3YbSjY0p7jnwykvZvL4fACiP/3oyMc6Nsp6G0KZ4KbTSVtHus2C2S2LespL2QO
dKmJ5n0LoiMEY7HziN7F4Trw2Rf0fmudL/loVUfq0KsGHqGY6eDCGnDpcTQ/6Ye8ySSbPpjH6iLB
rVoyllwL/ChtbzkP92dZZbvvGeOhTwL0RfNl3J1N6fpga5fGbSmu2dV7JEFQA+ecdh4TbxwKV0nF
iJrEF6UwGq70oTNHVmg2uGOx8a1paLHdyxaazVsk6yqWJGaHeFv9WC4P5QuNy7lwfzcuGyNfsNlP
zhasH8XC1IHGkwZXF00lXaBFAC4MpOL1tlPFrOQ+iXZCvmCEWNirFCniZGRdBR4xOtXv/dUjMLJO
RHZLjYnQZ1qaguUFyRZ3yijOegaIWCeRLPRnHeYrPtXIeYIYX4bYI/cYErLN+oYkGc213v0wBfsl
SIe61BDvhrkfrcEZwZsLnW7UACpbUO+E0if6Sjm8EY55QINWuYd1rOttmYGQ+OAxiIiVTKWyk+mC
ZsMxVkgRvAE4M4puR8MQxcILL+X9DplEb/PcxKSNtSw+kLXiKNs6LJFhFusb7oXulMlTwrKnl4jN
2KpossasK+3lC4WJ1yH0OdG6Lkn1FjWbr0Te/Tj+Z++TcZVzLj9nL2WjpsSXcMfW7dKX3zG9jU9v
dS1CBkuhqqhn85ZOh8Ggf3gLmIqOcWUayUE6tpx/qHx0/Ia+tZjdYBEstwkEL4F0BL1QOTkG8vPh
npPUl8r240ztyCkH3UlAuprqI1eZbftwiOAMM1gfklZemO2g/Z814z/sfSxBBnwtLR4pl0h552IZ
iHlTZuGgYKKIbZnPdneVOZpXaas/oTHrYTy31BLp7bwHKUSlXOANNBhprrgLaKAas+4Sz7jn6aQO
5uldeOGfor8cMUmhJ1T+HnrGHMa1MG3jdFePFil++8UMr4BrI/8/SG6BSIITQ24cNcyJILKdesbv
lfQf6In7dVN1/S1R22LgHsST14eHw8VrZh+0IB3o5F+zDsUUNc/GYeoFN+6mb9TOGnjqX4HtJOlU
r7g6vY4XMMZtH3ZQUIGUTjPjoVwRR8JYdX54aMSgfydMGhe3Ih6GAlUTE0ZCCC8cx9X3oOGHbICQ
9vLnVSpoXqXgpFaF/tR7Voz/Eeh1+YD0r7ks7b1uRVxNXzc3FxcjVJJ3n7EetMFRh+t+FFLYoO4M
t061pFXoPyhGRSRVN3GPn7EIxC6vlSavOqAVkFzhEYYycgj4NhlTohzxlxXdKgwpWbg3c8MipbSg
ygZgec4dE1wvJQuE4mEYt3JiRI3DnmumE4AolZzvkCp6mLpVttuDl34krrKL8t/vUEluSmXEXJbt
4IsQaMENokkNnQLK1YlhCOYR7KDFXMD2sqHv77KmOFBoouTETqnXEI5j4Ieg5DIYe4w2v336peSe
QIIOWxAp9Om/KpC6wRE+dpLhSU+xAUoBQSVLIIY6rke6dq17Rk29IhtjEZPj/wxUwss8NswvUl+/
52P0EJNt3yv5KvEtLRNPE8UVqR8pfUuZIHopeTyDBOdvj4ILfeh2lME4AtgrLFPc2BKNrrDAQ6rg
Nh/XVFOd65UqeV5acIPT/3UYpg1hXR/9B8WGVvJ4R+UDl323KDzS9/eBVaF+W22lc/OmtSSYQwNN
UtfcoIuSF3gTGd2wntZTqgDBHyQDthNoLpZxgY/3A5Rtg+wLqr1qOsmbtKVCQTRreKZqxAGOJO4u
MFOkCDK6FQ1CHup5k2VgZOJgHJIi85I8kgFMXWAML6opWe64cofykTrWF4QEMpMk4PScyYwNgpiB
TAeli+CXK4zkju3dIIDaGHQKUJSFe88grB2fKVmLcO3j1Pu2vU92Qcyom5X6K+W2buYtt38ULtW/
v3h5blY8F2znhOdtflcxk+70bXXAL+fMXQZxOw0BdHTBuFi/kF1ZgOVsmnTTZNjaJDBxsOttDTEx
4dHggPTwLXadtsDHkSnxcwHqmNBS8MfOeSnEhzg2fqdPhJ4tvnUgFrpx5gwOrgTVqpbQr9IMlWZn
rCJvZeAi1QTSa9Ez81XShRI2ZesN+0BbCMEY+TDAi4Y3DUtCPSxjQWFezdbIieaipvmdyRTRghVE
bTv9DmselL+wA8ZMQ/mNc9pKqBRomu2C6/8TUIpVh/ICrtjdtOxMjNDPEdGxI06aRUqprMPMFDBP
knTQKCG8Hds/Hi6diugLfvikR3fE6kIzA58QsmoZc4q3Vo0ZdsdznLGu5uh1okjhWO0OwMNm12UU
AymGX+QW2IIRWp7zJhr2egrfsMEeCa9spghI+d23sxmtTJKJNOGOcJkdF9W8YyQDKsN9kriy7z0W
BQbsuj2FaforqBHlQ0/2zZ9XjVhvxH+x4IhQM22J2bgAlgFMhfo4Iw2iRzyLDtsag9oc4fz7aa2w
S7H/tpsSNKRBKscxHE1QDL2MYg+30zlk9UrAyXo5PQCGWXnNOf2Znw1g6h7t3VeSypBh+X/Y/Zwo
V55FRJdvhKNzEpIEYOipPb5mfoPfLL4/AYh0TUhUL+q4uRZMFpO1Oa/Mmfds2vp/YOlyuVDxxZwk
u+SVspufU+/jajFw1bycFMcGEUjVL4aMD7vqmIRJz0Q62OYLx4Vhf/Kn8F2cbFAtuWL4vjHmdsfc
O4DyCsgd7D/Q2YADeOHxDh7XIMbvAzxutmsFd+IKmMotdK0t2EAvhx3dCMK3ee718ieHbZourA3+
JB5ON3QT8KvjeCTDr2eYfStssduFpPHemeAZ3MMx/rENTY9Pz74SXcikVemgm1eoE/2d97VgGURA
TbO8E8hFwM3/5XkDAaTPZWRT7TFQ+NGV436Qb/aZfDGs2mfiX8XzeRW+mWkwU9M5xJY9vScFJ4gW
J71i4wUeikp66CuGwVQ8afjLlUWSTTg94DU2FjXC6tS3JefgmBpUxdBnlYx5R5ftn24B4YgbP3/j
49UZz0MLuHJYZnjfC6UwXoah0j6OLkAqA8zqVzkG/HcEhZ7s5MnA2jkVctcVAAP0WhM+sPTdxGzC
9NdYNLJC4K0EfLs3mik9K3jq+6ktTy0Jrrtywc1dkXnt3YUyIUxu6laFI+ypI2O89k7vx1zaC95K
0j7lh4CtlOSXa0pNMpFFifWAhSeICemDoQUTV9kUXQoyOxJVBydjk7rB2VGAkh+601sMPv6iXMCA
o9y+cIE+hZAdmMwqMgs5/DrCdl9WVtI4un6twCqajijhUtjcFbwMJBHVuEfq6ZIxoF6gD5cWgpb1
+PVfbk/ffZDZAHPv1kwNSap/4wTgWlDeFrq+HF9hhUaQYTbMtOiSFNVNqMztqaxEgx9DQqZmO2Sd
ihHfX3YaU/3M9v9YYmAr1pxHgvsx84mX/m2vQX4InpIE2VsvbYekMyLFujDydtJF0zNP6pDPDG2A
ose8qcvDv3N9uMJAssS8IKEDYHzr2SaGDkXFdZuHrmuNl5IwJpul3eJVn45lCIruXo8S4+8Zw/AT
DFZXNWMIuVmjQji+rnkznegHFC9/MxWpDQyltHZmPmk1qnJ0WEwhF3Hkd/m0Xw+qlBYWJMQqpg+i
KHTEPmfL6+H7gVlAZK6B8xi9q+BmVzTHXVkkBzANTg9OwHJ/wJUptR3pT4IoLzmRssYzVKXQWUwc
j0ExKnK7RD8isbpsS+DPs/eXsgFGy7w14MJPbAEwTJnjs9+spr4GwAE8QTN31E6aHy/0WSfLpbZQ
df+ycBNLqla5VkoBJEoCUaXhKaIJHmRiq9vc0P8k4NIsCE7s86V+pSbstj2yVt3UauQjJOciDrfl
kKTMC9cS3Z1eOXWeECkxWM0N+twL2gHvjgMnJutrg3T5qMXerEgZEHIi7TX34bPno3EC0UEbeh2U
QLtd/XTohn7onEek6ZsA2OYa3fSRMVcB0jQxOddmri4OnxHCOT9JRVD1l2zRBQyL1i9C684U1F9F
lZ9ej1+Qa42qxT/ILTdkllmeJAtGy+Rc4wfTqQ9D7dFwP2iwoe0HncbFNiqLzXp7rjtpvjCRreJw
TqHoQTDM2OaGQdZNyXDKRzv/8gbJPMvC04Su6Elu6MAlZDGQYfN+pBXyT8k/3revTBwzWLxOuwpQ
TMfal/pxF2AzgvdCeiH52yJAjhB5wZb+sdSP2MqgZkFVSQRB4EmJvOsb1DrPSn7h+xSnE1zJF/12
9mqtRIOYYKdpGrbZGVDr/wpF9rTdS8lY/I8yk4OvnJGAnR4wGJXTJNmejeAOScVOLsekrZkZSWbG
N0vR23kQHODu94Cx1IUdGtVKyF4EtYSQ2n10QrtgB4LtZyI7sC4lutVtAv5kgqjUgaJZMWrixSsp
pJMNBuf+zgm7y0JgqB2bBLS9z9S2qhoIOO0nGS7eA9GzgDnYfyRukKahmIodmLj1sKiwt7RQiSVe
hBSjQ0DokWuW/krppafEYry5S1QrKoBmIRah61T/Jn8yp72c8bUHlqiKjj0RsOgrUs7k2q/9Hp/A
86CHr1lpYClEK5Rqtbx6wEnR7Muihb9z/ONS0adY2yeF6WWuFYKyYnNHBHc8b9ncSF4zlt+oSmJz
58s3jz/tg17jcwFsMZ4FF0H7b/SvIhcW0Kpe7BxPs4V+VYIUiuScreZKkw6UCgPR51Of7BVLEE3t
ck2rWhpgUbwIrqPhV+g36Idvx+p3JiNSSu9pQ9MgNz5h/tLWq+ZcoKT+yJOUmpDXyWPfYIrTCw9g
zXlbA7HSHRKcuuyJHq78paa1bE3ynG9+mnUT4rTSCBqztn3Lnd8ThWMYNazXJoVnqk96/ZD66wPR
uhSaXKCjz1JR4SNulCk5SWj8cT0OHuS72N56xJ1NT/nZDjxcsdVtWtiizeiqSz5DXI+mss7Dm5Qg
D0RmUmlZdr5DXs8A5cz+074Fn5R0tiqarTC3RBukqh5aOf+eKU9PQZdikgMZURjlJhrDX8lGTO/q
Zdb+QO6ZWdaUbUWnJe5o1hsIyUsWrXx2rvh0/JIr2Pnz8cVnwAI1bcPwRPvNVzDuTFCBwxHwqkw9
dNP962sAB75p/Kc7oL4TaOVaMCUcnAUr55GYxVe0pm3wfvzcKtwVNZsFHmOcxK8eBGt/yJ41Sjuj
HZmi0OXL/WJVCbvf14nZaN8Fyl4nGmbf5vNuvgx8+fBuDgQT494l7W5IsuzrqJNreg9osmIAC8Vq
3+m5lWfX6X6Syib8paxurmM60zMRwQFKrS1JNJE+PgrmQgwVWSN0CItw4Cgldm2JMiwJV7Zm42ai
fjhqu0uDMdpaGas+SebNmdJjYZs5alQz721LVZCU6zwgImRViUt6y6STwkG4wzqJtYBvWf+QdoMq
84GLJ1wy9eMgG9YHUBP5gspG2DxYg9lHWOaHUpTFnGH8WtNHmkNM+yaIf6AoMa/bB3t+gd7ZdEK7
omWPtPF7+5PIbdHI5LpjyQh6KXANGlQLp3RlWx/DW0IQtm4o6VbkMVap2Ip+EqdWceYVNEhSrBPS
Am7nUSzjuhkgHxJxne8oumGKfpEXmNjg6pPukhOPQqMia/Nxnk4vVU3DVPCnMTeBnV/1eqZo1iRV
spBR59BGcbkGyGXxs8C0L+21aBnP2qQDYToBJxP7IxACS+u3h3XhIaYOsdOxXxsxwJjphcDacc9c
bjol7+Hm3imHu+P69HGTkaVzbzJC/HbGAMTgmt4mmgQOyaz23m/yuIyrwLSM1ttXxsyTcf/O2+fZ
h5HMDcYW/Mygt/16vOswCwBgs00h/oHIaZtPiAy7KnSN9Uhe4374oW5MPaGpgAafhRKJ1T/ptqBg
6Hc5fjLWEvJC04+yUtV269Yh23qjlYUn5h3OJhPCgpNunE/F26k/kg78HtwiCxykErOr0IFTvCJT
rKXVCcDxKA+JHmstlZDFbnNelbxGu3/gojwbUIczZFsltiuRAjOtwxynsCyR0JYNMRsHsg9cliSD
H4aX3KAfZIX/KDA/gqo7G2iTQbhL4UhHfjtkcrLIZc+e8xMiWv+SqYl3r9TPkYkeC1RcVdzqh5uG
tlin+be9njC0pNjLygdxHTi3MDV4Ec2sB2P7QhkPrfue7J/KWISN+Rjjm8sXciogxoAncVzxGZNy
GoKuuxN+Jq7nyWASgh3Fld6Ea041SUvRB7ie4yn84fJ55M8CPD/+2KpDJMcnTllY5W+Nbf37l6+4
NhIAANHe/7DxR6nFr4fwY8ILJL8O0XGzk0PZ5rXJh4W7WugWED9bKPXV4Sos+tzaorsB2Bl8NBUv
8IGQGHB373nPpxc6G4gRRHIPy+PttHTy/rRoni0pfk4OOWODdL5avFmmbBry/R+PhVNXJiZvI5Ys
PqK0dpCsiC2KC64inrJskqilGC1gYJAwbD5mJOOWKi/CIFRnvJit4G3ZsrxgFSH6Ri/mZ/UFJi3p
5JCP1/D30yw6AS+c50YGw2Y2QHCXSA/XR2T53hXy1/GkoYh9VYmfej1uaQVvHAHaTWWQdu6qJJp9
+NWe/gjv29aLQ8AlkdGDiLVqLiLONGxFW4BYCsCedUbtLWmkeMlPPM1Zthf8MtIyJGrlV0I40Kyn
FIpk0IFNrHzeb0y9yrjxoVzaeFwIPhOAXA7qtsRMUMtLg7c0qa+8yBHiekavIxej6pqfzib8jEOB
/mRe1f3Nr4I/k3VJao2smYR7XhxVxdUadcBMpFU4VZ0Bw6/ROpmsIKcUEWVYERmP19p4QApAHi5h
/aCIGJwqNgiSjFoVa4annRd8FYZunzsqdTppvwbwi/tTtLWf9vU+aprGY+wyGz2Gz5Z5kbYwaASd
vtu2+yXOwh4QiOG4HPNXOrTZ+4UjLGEFYuw47mW9Un+b1foyoX3E02hRwxLr1jiyMAQeQdEvHx92
R0j4+dp6zwqybd4cxpAJk6/bu+C+mgWPETB3tckZ3G7qXw3mmnIKQsFi+XlZbp/1784sZ3HmZhXf
H9y1ew1tP/LtmYLKHGwnTqoTFh95Urm3SANVwYRTyr3dcQn1MPO3eo0KE07LJSsujprMaW0rFaMM
lgnaZOBmY6tkEK4f+JD/JQVHoc8eK3Q+h3LvefZ+OTBA9KetZlQr1/HloQU2jMsFI2dkV1tcJEtO
WrekpIfVCm5m5v61tet+10Nhx+F5ft0ybWjeDmHKhDLETehN+gvhYExfYfb1OzmBkjP0q0izT3EW
y69ql9jkEgy+zXnuNhEYuWTpvlCDTjMyuzhKmstgGwqQXGJmCfUsSC7cOt6WMnsmY5uvGbPuT2gi
BBRQPklr/d4to7tJDQkZDIFXg83xJPLgcLo5mQzLGGbfpIQTbTJ+K3xZxivlMwUJQF5SrdEZfGWj
nGqWZZZzQOtkTYV/5nGxulh3rVslw7I4FGzta45kBNVhrXgfLAXMbIl6ggBwZAxH/b9HlL/eSyVm
cAuD+TXqPqeQQrbCErqYlM6291yxf21cxmOuDWCEVpL8/Rjy4xC/CAplfr0UsA2o/9sz8+KVoksP
0P9+DOnyZm2QDjrQylTe9exKViYRn9WB4B/RAQHkG04f22DC8d7zfLdlljfjyCXZph8fqWsN2gs2
OmhUdovAweaeQRIUtPyVRdB4gsJIyqxQQV3sCV5SRqRLFPl9Vuk9ZF1U0VroTvRSrf7jzobQtBUD
TC9C6Holk0XLdYi9iaPHiXIhD0in3Ch913E/OWDPwH5XOC/23XuLQxm0yVm/uiIKXSM6MKU5p4XC
VkQetRUhi181UdENMIkwc/FG7Pbit3iAzx+8l6hg9/BOs0v1zQIPuF4SnSIPV9SJ8zj5jkQkrltG
QyZJmGIp8w71ZVg/KnqEHQRymDMKmRG9N6Ee+JUAryrQZZ+adieNyzDymSeWH4Hw+a85Jarsd0pQ
de5xKeAyw7HlpJD3oRrhsm/uad6iwsZU/8/Bd82UEH4Gs5DD2TsTgZLOt/lA08JuC7HKho8UDhmm
H/Gna3JiEM4zVq0EGfWInIfQ1R5PD5R48VHjI/yBP5EAorjAr0GGxuxZc9+2t+ieM56feKr0vXiS
Z1dlnH+D8ySW0OjIMi71S5UWp7cLHr+oiClxLyJRhjb2xdDPmATjM9HPETNECg9VdK9FRSSHCAZV
KivR885HGmbeyWdDULxRrblxPTEdv7qp2hWZnKrJYMROWDc0rcPV1vpO5lkb9TzfB1AeAhxIA6+K
0doUWLdaCiZkVYmibVakoYczdchFOHQZodXRcW28anyhypfsnLMU5xmhP5rujs9uQPBxU5KEQ6Oj
yoan+S98CkLQLvmfIaVRgAwr1WsfLzmYB1gAjYmHQ9KQUTP6HoZt6Sbk1llF+acqghknPARZXhKa
aBU9PcofskYQZQpZNIh1VZ/bl1f03d5CE6+XQSescUyalgZsBcDHvXwJLz7UNPokO8zQu/tSgOb9
2mLAaMoKGBoGbF4yrRKJ3u2VeeCIL6izRrXu1PegJS7cXxxbozhFSjDddb5YUTO659Xu04wLiQpY
FlaalylwhNq9/I2lFVqcpu9Wz4ABj6mIMs8E8zhwq1MMpeTBNy1Nm8LJeYMfC6OvPTBN3jabyyvH
FRam8/RK/OFRzxkLZ3eVJuVvPusPUNLmgeIXLbklgHqH/8tfODkqLFENSUKHeNmfxACDrsyXWNbV
7rzedu99eEzfKtSy7l3XhGfXbC1mKWO8xupT+4IkM5u5gvOC3oALofY4AN3Vvo2G436MiVaCqlqm
TnIT6G4Htafx0Q4fJ5Xids7/Fj0G0SwoCsN78gikcTSROuByWvCZQnN7IDv1U0xoIBzCbQFEtcL9
yPqM+ZZPPPezp31IAPXkon0mGBcsjWYPlEFOP28dovUxmSLDwCIYaNOXhb2ysQMCLwvt2sIwzJ6U
hKjmr9nqVPO37gaArRx8Q0q9lUwUEU9HVmlhBoXxoI5GfhoFg0JSZ3R99KwBCZ+YwiIISqKKHJGQ
zSJZgZOIwNc/bEZ0Z53SIY8YQeKSkW2Cg1QMpx8pOm2TE0/clCHFmWV/cIAWXSLOW7DHutlAqNhi
/7ou8z7T/DW5y+vyhuaWuWvoNRllBuNRn20LMZaNTFEjLMEts8QRX7HHpC5aAyIEpRq5BbZRro38
nH/BG4ydDM2WVPRQfg700eKat/yvoak0AX3wEA3L184+BiNGS1Pe/xNXkiP5Yy9dHr2OfcttHE7B
9j55kEVe+dQpaBvx9f04+h8hGG0hUMx28CD2FoVkn3gGyMtjJHTcxlC6XaQFt8Vy4xz6cwpg8jIm
BUsIyrZXJu6yi5IZlPnKm9T54jIlNoLVZsfxCLBmPRMRQ60VkpbydOr3Mhzr3pAF3ZL9YNx3qkKP
cB44gEhQ25yc0LI9x4wHVf9uV20GC7DYttYIDAVOJ18hRYFoAj2Pnbs8Gbp1Gslsj7wd2DRIkDRI
rZlGLhSWrP2PnJhhLOHBjI9UkVgxeBR5ezK224Z8RR2FU0sTmqGM8bhKyXKPRgoRDYurH5JzLpBA
5Wdcir1DC4yEqtDaEiRGniLwVzVm40TLwvM69X3qAO0VuxA51uUnzGEcVoQU6yT4u51r1uxTK5xN
L2lyYO8hwfVFioobDO+npLMs/XPewDknk8EMvqNYrcumu9Rm1OZ+5vf4sisXyW3p8o7MT9GqYvYF
yL9N/XKCDGQCJuAeNl6qA3eriszFPRJZY6mTgjCl+vfRkKiaJ7pAReMAMCTRiXjM0ltow7q5bzFG
xqedbfoQjpl63W+jNoABQeZy8aNlrHUqXtRIUaXPazZ2c1t6T2ukIo3POONEhqzLxEtyb4X3+h7C
qtYSjrnmIoZwN7pR4nS7SBUSXycFwuH9AUZk/RynpxhjSVPGoXnr/Qok71bQDk3nRPPdBwGQ9bxY
d90uP1c3njjRa9A6Cti5bWaesKcVPROYKNwQjWcvzMBlQh84nCnc+bBbCrUw2OwHC1Cq44UuhApj
f5evfMUqsVYPQlsez7kW9FT1aGc+6cpVGRvknMTwu2KLwcyf2buePM0ACeWqcs/sVu5mNKQLA4wL
R3tIWPCbIQybx5douZC28hJiSD+FrEKAI9ATpIlKBs5dfAZKgCNY6kcXaHUFZSspZR0mJHSCta/Y
8Qd043NCYLI2TdYTZEJavbI8SlFNfKoMDmfTLHHPaDh6bG2hDhVZEHpRyy37YdbajdwYnP0EPMiB
6Dmy3nQ2T55GST+/jXcQcYduq0A6CkoLZjX510cs5WTz8VcFpbGnsvfOOSQsi67YvO11YLhxp51t
Qbi8BGfCFWtejoYYm+FZtZPyJuZyRrQaqnJMHrzy7QIEjHmyjH+oQyYYaTjJqtcrAM1iUkIIlY6E
ukg9BHFBqQeQjw1CtmiMfsKUw11AMHVnxUc0HF4EG7xuwz0oq5k5yrAWi9KPa5iLvqEFKnOftY5v
SxK6TAbgufXT1wy+IOA9cqEN0dvFfmrNXi4Y6VkBdpxBTKQeo4fE95HUZSDeSB+Mn18R8Ie8826i
j2JvrtvC26nzKHNf5JvhmsRrEcC7/n34ATTw1ZftrchXeI28FTuVSJ+xgN0I1ykh7g/nKl729ybi
Aps20aSMnufnIuD/pcB3kf/mbhZNbbyLwf9CHKTRzxzlCgBWM5qonxssbSoJ4ANKqT/hAsNyZk8B
E/V+1lipvQls6ildd0eEeqcCVmaMtje4a12zCZrh1iPkkDFVjL+aU6CB35TsmrLFxKieba0nMr/1
hczXxslEZxB/SR4jnIYYQPhgsWaaHyvzZI0mhtSw+usHRKuXyjjWlDNwo8wM01SBT7/9KD2zwhqZ
YkMx5thSVtFVBOHTTqjRDo/nFRwooVEgScCOZf94cAbm17acsXackVRAoLL6Dic/MQNMO74LiH1i
Fp/GT/09UXS74SW3/qqwDxjW97R5SsSa4SlEqbI95exH7W0lB4OwsfH/krp+zWNkSXmZKqHQUknZ
rj/9OE2iLCSbFx+C6lzVJZ2FXp9vpW8a33qIi3fFQT+uxRPGE0nu8j3+VHVMK0pBjwqMVJafTasN
sbHs6vkArAHFgZHJ2ox+EKJCXrAO8QrzQy4RThWSTnRarMHUboK6ShSu73ey3gP+MR0sUNHefQTl
SqLQgwPXEqNC9uzl6ToBYAI2YNXyqRpI9B0oXlA8Xm0cWK+oKhrutHHu3sr00dJ4Oe4Thsd5dmX/
DlLWw2OLBBTHmJkJT3PgEs7FmmMSArOHhm6ndu9f3L+8tA2ixUeCENqSjOtdR1CRqygNH6k3+vmS
iudpzDAf0JLNEaQt93IMhsP+p+P0gYZiy/iqSBQfzA9XUliVbJED+PFDNV/CBIiiTPyWY6RnTfAr
A1NmRtTjDqsNrNW3OtR9MF6+4ZMNGAWVnm4oOzgg78cERbBNKFNLYtOoRxjzc+xvStfTfe5JXTb8
PCVlNjNOjT1n/S/P1LY1s2SKzyT+nCtB840rHtzmHemsnPa9b/2epaVX4Hc5m1nZPIzkz39zwXxm
wSOfMuaLGf0BN10KdSKwx9xCFb53XxgEHzNdMCy3c034GunwxF4Ctrawc2l+RnYEyr6eeiatjW5j
A7bcb5H2kqUdvQ2md7KimJGSHH6ED6j/IfedCUfFyADUcDtfiLSCdVf94TU5f6I/CsoxXWBfS2ql
KlvhpzhOOxDA1cjNiqAtSbfroEbKBwdljlfU54pLE1Pvrup344bwRsgaJNx9q8eRfq1dO3fuoirP
PN7bT1aTWfpeijrvghLDskJktCLRgTVAzheFisLeW5DQcEqqhBoA2CZjKxnv6c4T+KbR/ZU19cXr
wchqt+G5xk4iABZi7h3eOc0jA6Jryf/DtZGKnFdmCVnAjP0aWpFk2E0IF/3DAVEWtKVlmKKUrepB
SUrdqJoaRAKkgudtKm3NwZSi1pB5JQDpGHEk1ZOdyuh/kYLAXIpxgvH1UW7IG8ypm1aPs/deflhG
E3Ex9slFGsdLEeq9bztCYk+kJFmwR6utLIhXmNTqNHtu2xWPtYXyHNJWapMm1QbdZjoULOtIFvz3
QdCZnne+fXvu2HHyg2bIuktNW4Id7EgUq2/Ws0ZZYmhDzO1TLSKEz08DUpuePOJGYlyLaEOGBXzl
ZF8J5CW8tu8TAmFSjaVpwlgYyHvqBasxm3Bfk7/xhzdFYdzvMmGOyqLtwNa+NEw8aazSld9qU4qW
ohf9+PnvXJMDQMiW5H/ttYGhBfQRfO+5unjJEWVX8X9d8wXiI5aX/ECh6rKeIBIHOYKjIQsCOoXo
li/RV0r7+JGVq862Ej6fWbPjqIbNsuoDtHUO7YreE0aExEatX5l7I1LA5ZqbZn5wEFKCFwRUMeFY
TYXwXf/O8BVByb4MOJki0JYIu0zNdGiolvsT2qK3pOapiRFz1CK0vacAHXxX4AMKbiiMm85ZVcBN
hLlmc95KEY42Kmp4vpjS8aQB3tW9/hwESa4l6cXdKPC4isbi6kUMydCq2fu9vZUiEXld2Fy5xG7z
obuWIVriUaDolnFIr2vePUqkj47okUI7OcNAjJvpCVtDN5Y6C17enDrW5rjhZPeDuMfjNswK0GIM
wTBCxu5720DTcas+EGG/mO6YgydfcEVHEdbvDbyEFu1JWrghQr6QNcZMICkkxQz6oe0HdJRELkoe
7W0RCJjnThuxzlBSSZrcV8waSNIdr+gODhnXdHt3nl5++UUdN0FIHW7gATEvHPSnJdYWQFkDtP/1
8HCFzgbOW2eV8U9zZ2guZ0TvRcYyZKMP2MVeoAyhF1wBAb+yuRCagJ52QtAgGdsgRvubqGyrPo1P
FPTguJFN2C3CF+35brXQPsgE6NncW16vtlgTD5bVvBo0+2ef6k3IQmSnpl9xmM4mTX080HN8lgyp
UoRLqGvLHg2nL0sh2R7AJAxVSG53bk2L2Eme/fDZv6ppOKlYsZCxzPTRENsu1kTN8EWQ38XtTWhm
AS6js0ycuVCFDq9bSjC5W7U8AvrycHBgRndkCBtJZ3xZ8ew/xrMfUujYQTBQinfY+DwfWuKFxg52
q0tOMLw7pTUi393msXDh8nACCef+mM9++CCABoXatklp8EsrMO2tM/GiDOytCypLrgJfDoM68oke
kOkDwW9CZxdkwNvkCiuDzCHTyvQtNipLm06p739syVK9NjIrAUtTnxQClRFQxiCw5oMhOrlS7iD6
fxDgC2m4uZUmkDdXiZHwiJTORbBDFEvzO6RBeV5VyDalron3mqt2dmwukHKlpVTFqTYYnWs/e9Ok
bkVFnzT7vox2xHqHQzqPZ+v8oAH9AfAgnlsjnikDnoRmtt67M/VREsXPLZ+VuAKthSaF3wcs6NmI
CmXVZV5x7Xwc3OrtrZtK68oqPb0ndcBxyHrMGHKqN+7uvidS+SvBjbs3TQhXBvGoeoUFuMFShTxk
D+8Pwj/KHD7rQDGh2XYoU73ioxxd3CcgG7OwfYH81ARRTg+1hc2mgVZgcgJOR4/3aONyMj9MNezx
Th6qgKMwxYo1hrU5FsZ/El2C1xwacR38QyQhXuH2eFOogGi/3xSAIR80AsL9a0bvjbiMZaXduAXX
Hg0vp6P2Q1QVTrpvgHdcoNpD4BYhqsir926k4Xgl3eV571ZdH1k1g9iD6x84ryhLiakCMPiaWVPW
98Iy96mlZY/4jT5ZyGjp4fzNvx6PxUqbb+u5y1AclR+qZ0qWdrI9qefh+StNMDRStZtFcsIJ0Dse
usiuV25NBbisiFAuuKbzrJU1urRhtRbI1B85zUquxa4nAYTweLnbmFVWG/KU1RAX4H2LmmRKAvZu
pezcjaWUW++BpN5H0huU/kond1k7CSYG6kANOfaLOKLcXfqeCNu0961IluZt8RSWNkNj8FDNA0x5
sAUVwmYWiC0+xxKaMvqJPuiVRSrxoXys5n6uacI63Eq17zbCml3fbJYry9N1troJGSL9t2XVpOWs
l4F8vRYL/NFofve8qC8NxqgsrwnoBnHxxCzN9KwGIpBQju1PXFBX9EhgLftmkZXjD44exyYF8Dx6
DEANdO8n0qfV4y80/kUBWAla6ZYyiWKVTo1JiPMKSdKQ/VT2wAUpcF2bmOr4rwHNTrWhmf5C2gXw
yC4OTJS6hDOdezl/qHegEjQkkNFD2LWCp1nwi27QWJWhJOkoxSaxMkqwJwYCAkzM000OzStHgPeE
RLN9pY2Mj+bAREpmCaqjkrk9LPNWTiNS6s1R+LG6gFFyatTwYGDp+TBUf41K7z2oiV9BI8HcV9wU
s+APeex7196BvWD1AhfK4e8TmiPZ0AqJVa9yQFuynU0kUiycXq2sfN8hmVS+6AQFaO33Drc0CCFA
Rv5/fFVDVrsFlcV/5k5zdKmHWVrAwx7T/POa54ZXhyOLb0QJThLUbrrHMet611tBCtrY4PWSkN81
kKX/4kbm7V1XOr5+jTKGq9T9gMNne8d3CwPHFGNo1fZmapM8n2t7eplsW+D6PjWYu+g3NO2PTKe/
h8WJVAqQAj98FiFge2do3uy4KDghYzCDMgZkyAVBdHO+1J66NZUFOrfRKLZA1+1WFcU9bAGrTEwH
DZkDryN+1jAJoS6GNiE8DS1xHuHlHokN4EyF1ioB0Kaz16kDjp1DCrcIAVIXts3VbfO/ZLNgo2TV
QSp7kh+pQvYd29dQuqRDFdKF3fOy6L6m4SXXmc+mU1AOCfDNQvrSr5s0U/fTNy0i/rB8CbrhpFzb
8gy6CK9rmfrZ6GcA6/J0ZZZtHeyI5kwWjc8XkZ+wjufEBxQovKg/cYrwT8qT7oV8KQ3XSHEbwpj5
8tcD1fnCT+OOkEubn4LHGpawtshkhx8zjW9gHYau9Gr623BolP5+QPRFr4uvANMMIi7e0DzlpG85
2k5qyZaKtRMST/yOxEN9CveA5WneKI425i+3y7IDEynHlfLnBeE4rhQQfsBO7BpxoZEzzywIWnxK
1PwpebFvE8xDdqhi/SUaZiJEBcoblouUkyKpvjjobaHY3KvIBDuizwNxSWd5s5U/f1oxEQMe5pOD
KEFLEe0wqj+XC1yYmGgSN9EttYdo9hMmntvF8OS4JR/WeYS6Fa6C8HctbM18+Ju6rz/gLJdn36wO
/Gwe39OlAxWPJyURPCz8Xd9vDwIeYBGnKfr4xTL0jyMfN4bTHxd0IiH/mKxtwnvmA5jpqOaClV/L
I2VcnZwqgFUP9gjFvpZBjk+V/z3EU5dUzqsxdla1mvVVptkNldjxQdUNKdUyp6f81Zqtttmsiusv
5zh/nMBBLqDkFhzBQdi0flINsBs3unlUx5HZqiOd4X1nyt2RQQI3rI/n5raCOfYBxLF4nsADh2fu
54Cs7Rg7Yxg8Mw+eE673GdHEyMFxhH+d+Owj2D1rDjKAhLmxegHAlPgDCaVN+anZtd+4WtdRFXV1
Iiyk7yMZG0ix+OgkswMOmOsVAB+EhUQ2+BynBK1vvf2ltlxFWg6f436sxaNQofTll4EsQnlCsnew
dt4v86wXpbgziLYMWc6Jva4R5T3lg94ULeZWwTdCO2t6g2sV1VKtlOKkRBKQIJtJEEm4pa/Hecsd
cCtNsJjkD+CxyK/60CNqYqPBKsTbg3ipc1M8iNntpSgHKo34jclsLAeg8+Mk6k9jU95/+wu7tJG/
2XVB5IrFKLJVFUyH8InRXv9LLweRBnaiKlXTz6h6L//xtd1+JXzp0rEk/cf2Xsaf8zszc3BYAo55
U2xkHndq9GeLyROHP20Uh0kQa3c3dXgiICTDWlX+92rOlJVykftiKBW2PBAh27QkZam2E412LPbt
tGWvcr/vZHlB4u1iIsTsp4+gOyS5LrD3k4pgzTOoNMwiE85Uj01WUeL3QzTwM4gwpgddcfj8cBAV
QQDc2fjLRUaEW15fkfGTZ4aNtebWxGrmjtI9kE/LSbqTEMo9mfK9wY+dWKXfjpzQDtZ+u6QPxyhR
XXN+M2KQPCTC9izp6jv68JYj3aChUP7wPWxSP//yEqL51o2EFfwP8Zyf0mMf24ghkfbqZioLqspH
I6MuENE5FJ8nm9Fv8BPZ2Q5uVFL4SVdS6rqxhmwYgVYug+jDdFwBLJKLWfnoNxG9T10tGD1cxHKt
yNKxWPbJAjtHC917uGwACsQQAISYMqQLbZeV2/1TlF7ifQB2jtTO4+vhlWgeLCJLy5xSkFf1J5av
6GVr09pCHwQP84kDVUoMHhnJWhK5ON6HGRsNDNrwaOPq0VC6cLaO7SuayBVHUTJHHnwajhCJf71/
r6xEK7h7+hFlxmICFfxamnDQ2dJdrU7CpPoH29Lm43MQBiHlB8phddKSqIyOHTnx2Js+ukd6/cu3
/ijyO6BAgmGNgetrivVphzHCfd7LRcc8c0wNmemNnIkpTypIkCnA9Xjrj90FrPjt5LpXWiH1nwfI
dx9lOBuqsf2Ridqn/Td+O86EE87m1OeyxkhNh0JKmXMMHNGGEd5Vo6LKbPZOBbdxIDW1/qe3gUDq
tJhxq0n2xcVC6vKTAreZssxrY8eRMrR5XDN+X/Io+yFAHIoXufvdh20n9Uoh7xhqYf3LzDBhz8M0
ivTQSB4yL2jnmPXgiN82S6yh4bPZJseOIWY84YwkprGAhC/S26k/GzOqZ1A3rbOLIdLohQuwKnlz
ZfWB4YikPJKRfvwiQ7zdBGyDW0ngYHwd9HCT9h2UG/mUSSTI5I/YTPGPZiJskakJmT0JMW55MwrQ
bCOyVeC8U+FaK1LejuvvF0PLXOe6d/KcIdui11Iq15Q2CDOHQM1hQc4z398+v7zBWF85XeDgs1cN
qwS1psxaZccaKfGwB22UDqZi8tANfLDpliwRN4vNx82+1+jfccGc+T8yQMqTVXZ23F+S9YvdlxS7
7xZHKam4Xzl+SuPs3KdH4/svRVAcO2of2edabWjOD8Y2YRAnaIoMTmaBLom/d5wavZvQdSUgdZ9t
NAbUBEHkzEwu6W8hpkHDAg1hA0r6J8tmD5EnBni+wcJ6EXshn9QWBnVymaquDHRc0rtpZfQFjDPv
yBrRcNToNqylmErGN4spR/KN/2Im0z9Dai/M4oc7iWANOulBItjvh68rAfxO/LoKkrqwCz60piLb
JxcIckqJ6A7OvAPmsFp6kVPZbyc/KRhbH9Tw1n0h5hAuyUqhPBrAv/xiGsb/MHfwDhhMfwzsimNi
upbzZjA8IUEwI752zB7pYktyFEqyExq1EzS2Eq4YmxNMFURyG9D8tcpNzDGKHGxAjf6lt9KbKN2M
mHXSE8U+FPFju3CAq+7D40d2u6JqgjbuD4wrBPEguKlXzNcSBQsMTaAqo0Z/YBYQ/2MrEqxKsfDJ
7gKNfUFp6eQC7UKFPAIi2PIeKkgj2eYWrHe+tpoP0/aELWLmDhpvvA6ynMqWgvmORsW1kTxLzXeF
/ceWIpXdxz8nJ28hoGbFZUnasMgbqvETDQw48fA6fx5RNN98ZtlcTh0WKTuyGy74Kfbi4oYlyEJo
7Gbh1J3+1rXBvHrGbXZuri14yDFfPUMHqHyk8Pzc8w9Hpoml3IEddyue+fGA7QqwnNzP7w1vw0SL
0/bRpDzXbhnKT7NdoFrTLULDjMsmuZJpL2GaBpki0uuc0mG+L/SW1G2aTg82Xh6HmA/p/VagUvFU
5F08gDwJQOd3K+vEXbTbk3acK+ZnsuhmoiY0YQOtsUDbZj1CPcsLYmTNaGd+jUAbuvFizLmuH8ke
/KzDlT3nDRAPZgqT+rlg0fZkQMQ3I9gmCfu90uxiCIXyDFJaru1D/rDwulYqWfgBfch4cL/R8bXM
UtXzGrDP33e2TI22rNsOMjy/NqqEIa66cN5EOkQuvkqxGwQUqgM4vp57szT2uakE9MfkjY9qoMV+
gvUeexJ8abHTC2tdsOIQRIlnfSxsihF1VJaozV6Y5Xj+N1BlbicBza2Zh5ripfPA9ISN5XeOjubl
4MzTh9BzeRlm04/9LN9t5J6uhVNlatlv5qaR/VfKYNqtDn5n0AbhaKffK2fQdrBVtWJW/mk9TdoA
Xc/7WRcAlf4VXEgfeasX8nCu6QNiLWxRdBUtgqIi1+PygqToQIcYRSmCjyUKnPkXJlu1/UyCbgaN
VGHtexs0b8+D+fCpI/DR4bdxhm5pP8CZ1z66978raqZRuds2HrEkwJjLSRqjhxNgNOmx4re+9YjA
AiorJmUDj7JMn41jDuL7f5ifaIAkC50GLH1AKauN3EClGROFTHe2yvwePNOOFdWIggtT4BHyQDcl
fTTN/t+jDgufSNmLz7iL1+U0h3azb7P1hPAr5oMrj9pT3zcngABXq6cVoFPHxqPLMWaRuhA0797e
PWst3jPntWodjVU0An++m/ohVpGR+WxiweD+r+ZZDStYjxZqneMo21JRBqmmAffV8VTtRNBiRsYy
ypjtjHyZ/0VRxUFKCAIlucJd8MI7gqQnsl3GGJMiA5Q+d14mg2d3fz0C3AxjPrnvcTMXlenPJGQS
YyD2LWirExPG3Y2AS6QZl60JdegPOEd1HcvdeaddXGBAHirWMxQ5q7N0ruwbSqCEKXIfq23Rhjf/
+WZPMFHzw0136XAv5cGOvRGqQIxEuWD59961b/a4Spo3OJEPAuyOVRi0fvmZNFR2XbQXrGY/kEX2
uTRlfJwJZaxNmwwqReiN+buscsduJJuR0nq88MuxVMYeWirSmGwMmgI+xT51noFx6qlmiKOq2bki
tXFHFyV1KZP5ySGoXdT6b9qTMdnWY1udB2r37baF/RPBf6kgXpToGD8E65qRTaDlJbAqspXJjRQ5
u/pk0sOBNz1LlRXMTjjpMaaDb8z9N6pN6fmrWHODHM2isogVl5yo3HMCGEKNfM3+DPIFwA1sk7vP
46uMU2hkcGS6D1k+PD5b9LeNIKmzZmDezBFIpZ33xhqnljINIngpx4fIt1pLz35KiaE+xtq0tiQT
1ak0HfmmnthFjdu4Si7choe80yCsGNMVGG5uP7UXGA2SAoH51gOFJMKN9EF+B1jHLbSXq23mTsnV
4IED13pZV1NfrjSnDjAuijsmRjfzlyt066wEZBxVL7jL/VzWgcEKNNNf0LIZ9LQnMKSF+RdNyMgD
/ZoSEamAE6s4p2cNvAJQmkOVbgsrN95X5hD9apEnQs7aVLuOzCA5MtYg1M1dhFVRKbpw5SEl8fYP
Ff/Bdo4VQhOOG9+wkaFlPxleCHvt2rmp9Xbnj74L1sUQP8cx7fv10X0Sk80HI57GSRWNiQeIRiX3
sSb4IJmMabYx02DgnfxxOpZmrtSapmRTGExsNa0ZPx0UavEOSdngu5+v+9hhuTnM9hX+X5uM5O2L
lO6xAEZ6k1nxymTTX8kVyPtEWV4hLY3TXmQNcGicIiMm4KIMtFKj8Xca82GANG7X0/plH7nR5ZLw
KF4AzoUglu/VtUz53ZKLxighaydIK/flB4Wlt8wVJe6nzqGpcHk+/OndYg4zA9SUl+i7eEQ62xqp
9Y6dAF39MTwZjtX26mR5HhTWkXSw+d9Y4+B5V8J+ZiwIu4v72GRMwVgI6DnkV0qZc5I/c5LV3p2H
H79frNuR02m8OkdF+tvJkdz+TlONow2kzg7I7VTaSqbMH6zNQKE+zQcDGTQ0nIw/twxsZTSN7GlK
uxkvF+pek9PvHNns+OjahrQNEHKllvdGT51F7D7fNQx2IUJ6vWfp3JcYEMcTJBPpPK2JwdzmB/rA
W5imSIa+uHGUW4O4aaSUIp5djKpW3VS1cmbW30aDK12HBJ5VyBjx4nZo8LKGwIdEGBgTXPsdm4wY
+pe2ZNqcyTXRQ4O0ZBKY/HURxDr+FYRyHcZN6NsaLhGgZVwajeG9ojwvb9vMeIB8M7CqAOrbU32r
eWIWSDsumGfJpKRzFKIC+WSk+V8QrJKUI5W1IfFFVh0G96rM/wUo/DSUAqtFS93MFj1+la1l1Zia
fvuSSU143LlnHi38FP157Eb+oRN4INQvQPnaT/cMKen/wcjSoxitxCoSuovQgrf03khSvorJ53BA
ndZxDzbelqxId+lE6cqODoYpwdGjkUQjhzdxnzNWrxXA1jHgOYueie8S7QBwdjMvOIY12uOE6cLA
AoBgU9PgATcW9Y4hNjGN6bHF0RoFQSVLxj0oM09W0/VsRr4158D/ljTYxyWV+5C6w6q7vrWkfk6C
RJfT9tjf/5xURa0e5nEvntkeTIGW8rLkg8wumZpXqNNj3Fpqd2V0HI/5MJNPIfNsO0BQ8tsI/rTi
dBcid5olIunWhaVnXNEKiY2cfqtdR4XA6M/b9xboURfCjtTZ5JXxo2qoZXrrxEvaPSKAr6dsakIc
pURRQASu5Q2BpfvbAZfeAruaoR5lXbqmaUOkJpw0ybtybK6PE0G8D0e3Hwzvw5wh8CDPnF9+PZkx
jpE3RK0Ce1DwwN48rHfDphXhF0L23Mn9EgWYYfNUNgR7QfF90UcwQgwEPGCH9/SdW9MZVDFR30lK
DMsRDNR3svfKDP1+GFPaT+1PpIycVQ8Oo9YRAAkYMlNYBiK2Cd7rG60dAN4SZrjSTmmfz0njA6s8
M12HpXEVYEHN8fupGDraSv6yyGgBiaMr2F1DugWVp0/0552FOVwa+suCkQSMDn88bYMngogXxGgK
NiZiVpAfPTqJ1XEwTPVzmZ8HfGd1NS8LME/54iqnr2f9gLwSRHrT7s+ksygUSdUCRx1lM9yh6MdV
39lyTStJgwNdaNdMlYfDeMm3aeV3njw7Pqo7pbOOHvG2JccjUdPsK6AGCo+MBLwBTjm8u5iBJ8J1
+sD1PPaicL4lCa2Or+Eh+wXPbBzcvfmC2aIcX4bIdjDcngrtpgtI8QtSf4OlWT89g0AxvBlzB4Ao
dVcPXv2I50uEx0Xy6OkfySZqVb8ulDzH3OqTulwRca0xjND1mF2f0HSWzdO2djefBy58mprkjD8j
P7/TkiPqkchSP5/WJrBsla7ahY2Tzs3tdtswtOdchm3JxVICk1INnTZE3lJAJzPx5U1gbkNb6V3P
DW2fOA4hatkiV2+qQ7Khw2RmIk3zOH4UdXWzuskDRBYU+pdUg1C0THoZd2kjmYnerO4akZqgmbH3
pdR/Qnxwpb9Y1MxefVzcvbE4zMem8BcLvErVzY36RG5staLViMfI7A2KxNC90TDe06ECvFiBKk0h
1zbvaRQg7O1r46D6TJiMuWmSotxg7K3hDTcCXLcQFcgEY6VeEloLv/TLt0hDP7c9SHNh/q0ZBPVf
sF1/4KOGwwJqZeziZhf1ChkYOgeesqE5Nd1cw6mUiJZP3zwuRj40MHkWQeLuL0yNwAswRbdEBvox
q+9lswEVvV4ovhl2gRh0MTDVHHS/TFOgZhuRhjJD70leQtFsIFJSQ3rETK1VLdrWk01R6KCspAO5
v7dQ0LNwrWJvaFNZ5GNQex/oS3EFTUhL4PKsmSyQR4aDzWXiumE1WnUnQxFv4INRo6pzfoB/c0Bu
ucvPOWpL5kDbwacevehXsrQN/BbIUHAV/9QwCvIw46z5vwy7rw9CR5gBKtV+K23Vub6ttruDsxtj
JHYvHEeChn7QkJlZUY9DVQ2lYB1XKzCNA+MHCqOhrwaq7De56XUv8w2CxoJBdIW+YPZGs8uK2/34
plY4ROmKCznGf2MfjCYp2p07JVAu3PIpfLfk/qtQRjrrpb2O9lb5p1o7h/ZbUAghz9CFEG7rdPkc
DQiaDoJjmwLO7Qy7vpJ6SpPn0p7B6S+iRlxCseI9DFlRCjCIcljf+DI6PIO7oVhRH/OAhuU/Ir/p
j6VcEgRRGATBkhrUqknKuQK0YXUXsZ9/6zIKxF1/bj4WZngd8CjNFDl9OR4nyLxCAN4a2NUaBpAD
YXZZizif/ndqbk6xjYsQPgvpFFj3oT4o3lkhusHBxeN6RMY9QfneQtM1leab7XhIuFU5CxyjCpe0
wY5mT/HI+bMkyzcbxkc5/TxRk4fp4d9Y73Ha70Py/Xv2INpfi5JugK+6uDU/JIBr2qtPdC/jWNfQ
soaxbL6CWY+/8rEk5z2hPScA4VO5l2daGBTTHBrYfirvcZ6wM/7SnEbUSSaSy0mm3+omAaBK4d2i
s0+YFxLCH76xiI4rUbfRlqFOiQO0oiWcrnBuuT2G/f0vWS/XbHWS8bwNjtNubUx2ELESyO5q1DDt
x0Q+Co3dNfgTCTJEuYNYUp9cp/m35Ps4FpOlUoYJtZn4Voiuiy6Ghl5gh3ZsDzMNkXsT3YIY9pC9
BGqOef4cuRXfroX2jX8jwg0qD0qRFlYQUN2qq6Swrf54KiyeDcmNTeFGjFXXXv2b+YRtEQpxGW3P
Ug4CjWgSJu72Bm/8Lk6m2HRSRv2C7oQctleiGv+2XzremzesdNuHwbETtoewIZG83vxNwjOqts3W
Y0/ZTEdENSEPumHKEkF/jH9b4MaqTAXLwqjjxAOrxaIIMMoZCtp6UeU5Qjv5XZCnCBnV51a4PsUC
yD5BeGTbiUWB29gAYtBiNDq1zO2k5v6n45M8sbRs1SFGk+2IPnmA0ZtB3ydafofU3FfMVUe65xWo
zyVxxhOzUREiGu3apaP6R36wBFT4Wfak0JaqpyZXlcrzlHqy29L6tpeHJH4BwLDzXyO/SfY5jFSX
rkPfJi3aVvxXxjFDEMxQHxQsilNexIcflCVz2D5L4msFFRhbnXJ0ITWLmsCbg5HKFz+AnnPoD+Xp
85NS9vxYBjorz0TOGnuao3ohZg3fRkECzCmThm3dvmZwIF7OB2yz5M/8rpum9xQrxzojcvhvbSD7
WRIBV9UpHG+IzKHTOrctQWQ19hocgMlW0kfWjrFhd87FBHpX7wl6WlpwWW5qvZjKEc5xGUtQgomQ
EEx3a59PWNLcW8L3OyCdWLza4zLwZMlHn/bQLfoybi92lPQ/nF50mV3WXQxr5D2U60/pwweaBz4D
48QjqTOYgm0sB96qcN+POGW8ncnuym1kBsSDysu0a7Qfe8Jvg5nNTjEg31OPSd6RNS69cBPNpBS3
GrkcyP2MWD0ohHtPkwItMNn0c6yK3PlHK0L2wNPtH3rsTCqfxon7BZ7uVmnl3KPLlCnaYi9p2FkS
YCGesygceoPOuirXYG3n27snHzDdKJiJhPqEsxa9mgmPXO20zFsPpiGIePUqtwS+0jPRMuJQqMOL
sLjDzFTsEQyMKbwyXhbIEry5OtHK1pYEz1FEIfaauXrUPaMNawl2HhizZDwRRMPPh+tQ5iyKXDZw
VDae1QnmwxUXn0/nzvZmj+vdlUruTQn+2gJR9LHzWdM+9IA3Q7DmdoW9a7cpDnA9CI8iXMMi+Zqn
wwMvzJ4k7Hg2504aTHsdTwXqZT3PpHm6Bm+Z4Rxlxe46l1oYiNn6XmGr2vWUbovfV0LY7NfyRGQq
fmXyephoF+bVBaDYFEwwN8HoVF+n8Kb72jo4HnM1PQwkkQmeqyPn9wxb33/yk7oRnVPn+BkmsL5R
w9lLwCHOnp6VVkfUmbkMccpOzNPq90jTMgRdgdEd2LmAspe1TiYx6vOupJe1SLI4RsixDLlGsNhX
o42ksu1eJbB+eLDPXSfaQNSBHi3mQDUFGxjQuHqKCvaBJn7mRCEaPPoBLbovfQY1ggf67QdwYXF+
KdUP11vnC90gxAQYkAAPRII3QaDv3etwrkMEmwddukBOwiOKehq0WMZsYWIAHhMCYsNhT7uG/kqC
4IOIvMwEtc9Fro4C/5Vta5ic7l15/+7MPzwpGxVCtPhcPhLjdcZJ9vHliiy47Rp5WEMGRByr0gIZ
HQuJcYrLx0sGrakLw7xasPcS6zCa7aPAuaxxBOv87Xaz2BRATdcOze9NhSDri2wfgRteOuQgnnCN
vPFZkcio8jRGehmELRsS6ZQdgpqpJ27aYpwb68NNXmAMrtrkmh4nxDK7Pz6gMvORhTxzUMHwJyFB
g9yGrPxqcf2WnhfduoodUUezpnW4rcHa3zHknrGW4V9bIZ0FxgnLNwNapnQC7igh45HDEyJAt231
TVjnMAiuDsld/tyhwDylaq+GYJTMLb1SOmZJJQ48Zf14JziH5pnuPMNVnWHFCP3evFHb1zljzKln
pPTruQLnmqj/D8vQ9KfPBt1mucOF0uG5wxuHyivruEnX/Qp6pjDn0YEUQUVTXm5RmMw61qxV9vnO
wqWlizwLJWxZFhJOrhSyP5tYNtx2xsFAKauWrQIK9W3J10fFd+EVaQaMWQ6iKlsh/nQM3d2m+M5t
QYBwwi3CUTSoZB/qwaQXc06vip0+RhEBd2wq8F1q7vJZmakfkHluR/6LZrXmW4cho9ZpsI3uZLiy
cb6XVb93Av5qYuGVOX5ZZksVJskz6jQJ/XYxQkQdjWnJ1eLwurPc4wWzPTRJN2ntprwVA5HBTYtc
jqeQyVoiMPrhr62iZf39TkuymzHQ4D12G01uMHJ2+VhpsS+hQN58OtMVDfXG6tzdGZ6zBvUyIWS9
FIIQP3lIqDGtAlzt5b3b7LmLlFFalbOKW3SMdpZEACrmNAS7q5dz+CjSWrDkg+jpjPf48YQ6ETyc
nCBEVdRbhLBJ/jwpwu8WRn6XHcN+qPWHmqgOzTiBsdrQKh5ado1YWT9bSlqR/tK81QOeI3B6o+s9
9sy2XnfcjMl3nhYEp9VWaJqoHUCZyBoiyHsM4OkJDfGIbgrmtgVP+KZ47sAloCO92fIN1aMQpWt4
MIzazUwoF4wvCekwV6TydPUnylj03KdSz9L7TbeTxpj54mWeGYnvADimOc0u8zKqhA4GXwB12L/u
Qco6cx9bTcyCtgdjfDr8mkfxKOTI2SMl5HDgXauRgZEpUaNSe1PBsw44T7E2IKwnqZVlYNiUTghf
6QJmb1VxOCdK24J0ijqWw1DqLT+zdQ1VMzRHE/N8LKz/NgFh46eAsQ3OTpQxYd1mPQBexzdBbBff
40LMpILjUNiq4BTuhoC/CK+wy6LmB+xAokZUYfJ4rLwU8t9PYpyS4hRO3n4A7+9lQbSXEqdO7CE7
K9Y+Bhxg0+yxk17g/9tPzdXvyucakaoP7K97dzOstsO6oO0yJv4ZYLlvnfY/cCvgNESKosxKqiCx
odG5WrFeGB2x2upVH2w9RqRihW6GvcTW3aoe8mi+8RouyxpBlFoDRuCJVfKy1bXHvU8XnS5/K88L
K1//v2IlxfuD7KzhrslnZqk4HEisQ5el7tF0uDqUCcprIepuOwaa69a6iTMnZCkbYAQo6RfevueE
ZPU5wjrGfgYKweTcIg/rFj0yAoZuvUwB16DQPxQYhJftbn4FReg2rcUCAsXe8MRKpbCIpve+f91O
05qSXxKqnWCR3NnuSC2KJHHWYeTAyVJPy0D147b8V1mlmjSZXPbyP0C4kU565oY3gu6KuaPBUgoF
+VnMI+PgkfuCpFQ8UKLbcUwRWh45GDfodGAT6CLmgn2sfpkilpvxgyDAIT5EE1Lbxu1lk+Zdm2Zn
lh1y4YZVNvelPX5dI5wDNQOICWdcG4RJQEKCfSPeeBpC1tW/eKkO4XXTUGKWXEzDUP1e7E+rYK8H
RqQowKMVbz6gg+fYPXwLJisc53+ntabC3ROA5+O4gYYLpfi8AqW5XRmQwZpRJ4RVxX7RbaK2W1HX
Kmo7aeIDMwy1oupT7OHyL4ZVTVwm/HVzSfuXsftqh5R7JidbgZZJfS93gsa3usQbw9amHBFQ0bo5
ok9KGeBKIP2I/ca3Jj7uv1eW36y/luiUCl8GynEMyJ4sgW0JpWDOLjhmoMUqAewmXr/4iG0Mqn86
KiUD7VTcjEG1Nqh4MT9g+A2r8KYaPTxsZ57Kw0JxQp7AO7z+YfqT0bTtgsLiiE6jgQmugiag9YAe
TcUa6MD/2397D5KuhnLFgknJ7WciLdtTtMzHWycmy3YQ31+K03EMo55UjYkR3UxhsSPljZ22Ap1o
hma6BUlOW6AGLA+hMg/AsXwyOL/hGVT6HMr8llKCYylsAvSLDaapshJZ8PrXzl/Ec3hmVlmQi8HM
r34Y2e6gy/JKCpy6kTyy6nIydBH3+C+7mh1p23mavZXANAb56+wXC7xMlSB5MmekkWoAmXywAiJY
Y9jEf+BfLfPfaL+SJkMgHVQOxbromzhBJ8K+0cAYtqH5ehy0RBYvHXOdxR3Qf4mz3KWQrW23fpUe
eHON68MBGDX2DNVjPoKXizaCd6e7JOPQC0R1wIH60U5dFiDjPdB8HmELVF+KlZ5hMNSFSXtvE/v3
Xchfu+gApsizGPRrZjouBnanKI9pBB1jNQU4++QMPPVAvo9m/dkTrCfmzs+H0GFs8kwraPi8pkij
l1YUGXgl8mlH3PUZvs34VFMGetobKvXhmU8UuxyNhsTGe3HM1l9NkPB5DPFl0BuzrdVXOjfvrobh
UNIuT7TszI36AQ6OoljtODrp32y0Vs4heaYVdai27mTOScji9N2Brm7WU7ml/vci0FdAFOoazKbo
TfIP8mxf5AE/O4ht7BH2ZaSVzstlMu9y9W45Yxr9F4IvJRzNt2V6UW2St0J02VYkYffRDGtUNjxT
AS8BTEXmtPJ5Es2u1m7mJwTiv4ZlRqXauTt5+cb+4s3wxjah+M8mZbxo2XNQPAJ6/KNXcrXDRiuJ
Ac97jesBAEUpHdgthbN1sF3f5RQFkzJ0S7Q0JboCGWDC/kKI8GMVeupkUy8gipdUft5SeRcM7ANo
/4hQ68nDJcJdZMNwQjF1wWU36uuK5T5rwYu+WIcCfrIHYFb1gJZLgpvZ2QLXW9Z8sEBZNl3Kb87Q
r8RUeFCB+frQrCme04FTmNNg7o8XHfPl6T0ifwZZfb388vMVVINvglMLF3gzlLOTJ/5HqZDlEHg0
VVNGJylbUlcX4xxtE7I4Lpw1/t7EXPIhSsYmiC7Ym/8tG0psImn0V13Ymc0iCUtFXzjzVp2RIvyz
I1hF1W9LEJdt4YnWGspnHQHLCZXlDRDxzVAbafnzKAscMXn9vJHctxtheIa7Sr3FQKmmu37RD43R
85s+p8I9xmtwo4y6RuERQPxx4ysY9j47rQ/wzJ1powkO0JxdCMOZGCnzJq+j6Sj8UAxjthkcCcNE
foXz03XOjfQ1XU2b5RmnLkAy1Sqt67W9lC3TabLIDrQCaM5WaGRWxUwn7cVnQ1Kupx2vCUxmG4z/
MA0q1zFbO/MOPWYTQ9sLx1iBl6/k8l8CZzQTVIBvQ3q+X5zaP2t1RU+65skZ/28qKboRAomcGg84
06MP95w8Mo8yfCFIeif13gmHyY22jyqC77zHavE2wRfDzq/YKkIcFe7nxdiCFwQ/BaI2ii/b7Jjn
s83lI718orCJptU4GvELQJAyh0e5MoXzjvGcUZJpnpr2fwxQM60xLDoMwhu3R2XtFUi14UPToSC2
yoTN7stpZded2wMzfHE0U6tcrsHabhpl3tXJG8I4D4qMcfeiiPjWMYYF9LeJTfINvVVb6bYTsS0R
XftyWq5MZnyFeDdL9Jc56RSsAKEGR5SuDan779H3mjgGBnyVqPawPuQ3zvNkcwxvcCLALihvv38d
5+kvPKF3lqcWcJIFfrCt94tyn/bz44ZjVrscQ0LsRElHAmbuI5YidZ/gnl4dpFKXSO4CGH1nY8U1
J+bE1IkHmdr4srrFgUtoppu5irukUgzBmSXeNVVSJyATJO3AXZIHOsC7bSNytJ5t7TJuy90MD/tx
zdnZEtUV3s8OcOy/s69Pa32mu7Mvlc8r2LN1Ixrn4MX0jIJk/tzdMXHcKvA3I3G0ZhMBgnvAMEPe
F2WIXVALezQfoASto3YlsbRpoIZT1STBssqlLI8P9EeD2zFgz3b7YZDRRD1292YSlinbM0M74jwD
1GVSkr0Mg1Vk/MGsE4z4HmFCr4gAfOk+VmesvQcrGbAAuzjCLnZPhHqeh/Sz7fhSauCd6V3HHdtW
EDgKW4iEjIyNgJ4ufbLXYXWG1HQQ3lkfDK45JzY7U266uv444S2Wwy2charqwAjgTLyuPIa+3mlR
B19MQa4ZRcw40R6W9hC/HDpMbuscy/iQYD4FQYl77YnyQFQqBxSwOX0xhWZT3WbrqGLMEtzabTXl
Wc2cpPQvO+72sV7TOrn8nctLAVzFbwnb9zIsyFkOTrZuNQlAvDquF58Xh1fYusZkj+0aQCBv3hAL
fUUZ8FwlGJM1WnjQR34j7N5Zb+9doHMdyUbUzTMMC8voU1+aWtUE/KT3iQy443GQdRRvB5XlGaU8
AsWvDfhJ0Wmz/6W0/viS+SdM9QFNXUAdfbDCnK+DWnJReBvgsL3hXba3aNi85p5tHEoFbF2dgaNr
JGWyG2g/QXzevl1kVaXzhzHkBhYKlVFsg4gmL0MkolvAckxgcay/vp4ZFLC1EkNZQBwyUekJhTiq
JHgZHF8fmNWtTYCDzu0zfjbdKJkvdqOC5FPH8F3mwyPv5nI9uVMtCBxC9T2p2ROM8jW1qUs+8pKA
AO/26hAUjqGf5R6uA05EajYlamJhjj/oswbIHp2qumUDl64tatBaQKioIBdxoRG+uY36gQBe6j18
cmVuqpcFKe1eEB0gNlbeQHqyC2x8EICaZQlkYDguKV6Bcya9siwR/DCagnLRV/gylLQPP2d+1DuQ
32ISmBZi9Cy+SoyenyWSfPAWlugbHD5CPMxVdIT8tHuDxlTbz0G8rv0eO/8BTHINFmFBCNBCd9MR
KeneYAf924q2LCRMYN4U4Rdb75jvN5KhqsiarqMfoULOyBUyIJ9YizPMpENo6xCzWsq0hIzZf1zq
nFUKE8SFHZh3rLOc+PfmFDrIc9ALOscqvP102Uk3Uml0ox8pzkwTn3EoFw101AlUsDG1YIrZfiuh
Dltz2Xf8KxBUDgmMaBW9wNGp0m3McRAIbPJleVmxO/hxclhnbx8FB4SV1gccWopCszHSo41IscGI
k4TITm2ZiOc+LiaDZ0Tovx6nfbogkSiFA0xO0WqRKDsOcnt0mClOyFIsGApWqbVAb9xpcZEawL3R
Vk0cGRSePBIvoX4bCJBjx8Eh563znWIiar1W3VUZ0oVs7PoE0TGBms9qV9x6WDWcmv0YZaN3EFOr
qLJkW07ksQZGrADZgY2MXWvMWGFnabM8/J+CaZiT8aDea3+8Ms8+j1QNjMzzgrA3rm+cGSggU5oa
eBh+ZzIAl49gmTtVyXDADA6DHf3qeu/YHTd27Cf1YJdEPEfEAQvmiq7fzbBsWL01Oiw8FWm3Hl0A
lzrUyhCPYGp/7h5OIyrNWoiVN5n2gujCWjfXiY5WM1xD9MXoqTWwvWlQo7/25FB6ogavTBPyDyxd
rifdrSkAHT7/9wArjFSibc2D+piqTV4mq4d7rxm8/F7UCPBkdhLcCbUD0g3H21R+gKCVn5yNkvOl
gMIRu6guyZUoL1qlxUCblM7LJYTqOnqlee9amdfMqLSCJYya6yriBCRpza5pWTltdATHk8y5/tDh
BT/YN9IxXE2LN0nhZiQSj0TmYvy6VcWpA2M9aUfBjODEA/Ul54ASrElSu7qQIk5neXXhvmJUT4Pp
48WPNpEK7Ug2XzQ5QDR3aCzqL0ld/IkSaDnBb0iNDB/EDKdF85PTiB4WdsV+0m/trDsNqNyrl0H+
KqD9IXifWL79SA41OA4wqXL8qAaSqXXETQbVW3TJt2MgwJwS1sFPkz5vQHdDrtnIhEukY64whaAp
ft+qi9gzeCGjRUhrTK/qXtp5xd/tAmEioN8WihDY81KjV1NWX0pi0jpJmOIwXH0ils9+uv1AbwXU
a3aZjaNA88KrZJdeHNO0WTZ9K4QCCUYFzRqPGkLWg6Cm8qmnzS79IpGhL1ZPXBn8tcoFKMiHfgWw
koQ6sz5soVnEmqILKZS6yk0iRRsiwgk9zlOGi4ywL/vvf7PZlZQ4Xr15r8EbQ0AOjjgzBBsxRIQF
vL0a+pT6fTZuggPxCHQM1x/Smmj72lfdahP/v/VkrS7IuKKW0wwQIHTL+xRwsLn19TYy2PVo16iX
Tm9UwtwIt2o4aei7xzSgwaHY0dqR8A0RADEYRK9gq6RjFDl0TDCsv+WM5sNla/+wUz++pbI2rPqh
0MkZnEZ+pi5IQ5IpQIX9s4Ur9R7mBmTsKrZaIl94poPAin+TCJqEUcCBLMkNYst23/tKThdYYZyy
BHXy3gjsQilIGAMzTiwxzsoO6NGzmFydcaxRxa82/+iJ6tAYfW4wH8sYthX3QNLr65naCPE/0sP+
QPvdqkMGx3anOg23jyaYB6zoRFMA/HUNA6BOsU0+ouH5oz/N8tSMSE5aNGWaEWZZ3UjTAV/dMv0H
vVimtW97+T9btxYNNlPi0j+PTXocgMX9TTn4F5tcBgnUoNUdtLJNbWtXLlxYBBp9SdxZuzm1QEOR
dyzmF01c/u0TDpJU+dBm7a2E7nXzHO1tYPLlKB+7rls/h/GfeT1oKP57qgSWjvR0/eJUzOdKdZb8
z2Zkkcw+eDDHKayNjY0eUn4c6CmLhEkXgxTgsHl+xof/bJRmEvqGK/iM6wfatZ1l938SuNxQc2E1
LMfDH5McOQRAvucPGeUO4boLTNm/Uv4G2MCIDz07rrQZkSjnEhqP1KcKJDeMdige7AIQb9dQRbSH
EJcvyklzJm8e0k8VH9AEgirirJDtKhhLkznHHl/r10+TTgrbId3fqOlhnX+ePFi5T27JlZixJ/Kf
wPOK6Z9QDmzemHURNE+C9ShIVxakee+DmtE6CjBvNw4qPg3ohbGz06SNZ0AAglebWQcNwuA3FW0r
Lj7wEDtaRplfnp299icGIU80H1OAm8Bmq0dr02BgyGW4FYCpebHMDPRC/M+j2fzE7IAZKi8jJRzt
jo9BKZTgXwCYcygwF940CFYJJMx58Ju6tZXFMY64oLs+WLlr5ZvHm5sXsFh2qMPCKJ/CVbgk2A0s
nzAT1jhoWyjFTUvZ976XAs+u/KS6QJrxhxBlTfcwUxLXw46UrY5adsyOA+s9qKVkXXQUlltrTJKO
V8d7e1zvuccPPbXCFrSsxKNjEmsNrhsz6xU+iEoEIvbxVhUvcb+e0lReLZ+yOWUruLYFTPVJUBVF
0xtR0vl/O2oAeoNrXulXCk66xRtrXqbEvivb4NsN9L+n1vB6o71gKobcLK3re5H4hwKa0r1UZhIN
rRrET/EBWIi/myCU4txdjWLBtebwcMoNpPVtL6eKq7cFQi+ub+F+WkQ344v5h2kJYHA3gOAjN+DJ
JBSZjhg9+9oE+fcIvG81HufYiHsYkz8iv1fu3pTKNL1mUscIaYFtqLRRy36Gy20+rwEpcqWYl3XU
UmRzFvFCkotkit/ahEUOXXwuF/XXK9lGBGnhPOD9N35xOk9cuWxRZGWj5OwUuatQ6v/JLEffvdnN
k8l386iDbhKZzPwYwFA5aGMb0U1rmegSHbF28bpFX9KsCqHigOb9IaMArl6z/gsCX1oCEaWJuM0l
7eNCINvVNIyk+LiziZHbG6zLm2vWZxjxJayUq33ApHgUbQ8NxcBL7uDavu7LDeFzsPQhLAb4ZNFK
TqVN2I/JdqANIO2kXg6+Wl3kZZmWZb4uqNhdX+LA7o1bftTyMvxxUPK7XOBVma9YLJ5ddmi8gk2H
hV4Ehil3nMidxTgXl6A5n+pNWCsBt7LCsX/Df+HVo2jArybMsGvB5u/uRi4FwVPYBjB16p9eFdmr
74uwQnGmaagtgCdlI7T/KPaan6Vu7IxACsadm52w/CjNa/rnGGx1TVDrmsjSs+NjP1RAU9Fj2dJ0
qaF7kzqajYazpFQVgEf+zOeyibORMARmwgIaILjxrNDdamWLt2Rjo1pSNDikeE5ZQZAymeDJGqbf
XNQKS4KUlYqO+upR7HHzIGvYBEFRRrnEgiIBDmr73UDAt88anFf6uM2Ke/nLyGT7QWPsHr4uzmLG
WMYoQbZcNeW7+WxLztlOsUUTjgL8m3bHtvSNH7XNI36hcfuTHuGSeW0Rj6qlVvvoyJE5GZq9ys/E
VLumju6usC12rppMSClfCxwMTXw4RitsnsMIIk0vxiKQZaLxdV7gTK8HRrLSjfHT3pZPUEjK1lXA
rGT9K3tCG7+ViMurpO9+j18Itq+NG07E6GOs3BoFinvhEke5csK/Q6mnd4HpCS5mfOUEwZKkkba+
mtCkiTUnmajGf9EMEx4s5e6BWNZUcJQ2CVzeIRZEshbWfp/241JXik2OltC0lcPuiJmcSG7GDKAl
eono3vtht4iF1RCW+hnTk8IBkGyL7Et2L9MKGoGCLWVX6Tr0dboPkQWWEFEF/GBc3FJTMoVf9QGl
1MKxsnAJzRVOOe5tvtXUkJIdqP16JncrtNnRiS1P1Yc9f8nyXtZZMLg8teiIoVnlSpmkVFqt4LLM
GINSlHBQMZIK2dkdnjnuBkzfXwTh1AKCm2vEwcjry1ecsgeNVzw1XMwNOgcTn1FleGYDLDk0w/Gh
/BHDuojzzh4iSnUvZJOoCJd31JhEtwfQXrNKUrbgdZjtKWZhVK6j9kpOHpan+U94zyzUZGblaXvS
iLAWnof5YJwOs0Tj4xx87fctNq7nG1PMy14gJfYMIfGrEwyC4DrIh+LYTwf6Dgvp5uM1Z4ApoDvM
2hPw1+s0hvvULF7Uri97ciK7Jxp7HIwPWcy5tRy+fkEoa1a1u3zZbKH2tP7tiGfsKOTRLkO/vrV3
nAtdUk+C3c5FqwNWbmnweZLG10qHBnpm/INpGJQcJbCbcoXunyaPqjLC5LXUOD1atBnD8u+xA4b9
iq/y/vN/AnxfKaGtvWZb64FvnXpCzRLDx2gxHtnKHbtyv6pHcd2+49syc86zJQVpDlHop37FKEfU
NduRBuJGfus87AlLHC7E7UfzgSIW0U0yaPYOOa90ageovYwE7Ym+Gorjpv+7UEYOEWUMU/3gUaYJ
ZsyUfwuOUfIFB1wxIVnQzz6xrhvj0B71kSKGe+fSqSO9m7ECm193CVg0R5BOKNxr8/hObnu7UPcW
ZUzY5tQB6EAohuQnu65/xWiauzrQ0uA4RAc3PoRWQyz8pfB6MUwioL8LBvSe72SVur0nOiz7F2AY
f0WSW/k9EF5YFGW0NpPgciYvq6dd/fxdcDFI6QlmATvLOsU8XVmvdZRBnHSNwNi2MMK4gD6b3Xu1
bhVRN4rLRA4Z+KqQKgSZS8DPYWYGc/xvGHRVvQopQY9/5tZBxX0xA9us7G4DTk/nMLpraX8a4psl
rI9uj/F84tn7W2Lqb4bkpK2eKSbVkd+icLTdIbRSqUOpX0xiph/0B2XjTZ6VYmIShlSRPoQ1dGKq
B0iQHvJvTpueFN0ngOJ4TjZH7N049nPd1294ZJb1gPbf/FZL9GIa6XDCDQbE27SXqVubB3V2IoXI
ytw1XYWTsmsRQ/4uSRqbo5mJxexQetVCUjl+dlNFLTf7wz+jMqY1SZbbIFiB8hCnG78SUfVtdW52
GKgF6ds+AlHTOhDVLKcsgKU3SQhx8dImZCFNtR0fx7DJWim3zZMYrzBQoSRATTaFYmpf1dyfkY0C
YSovRJZIvIBmHFSKcIvFULKVeAv99hrX1xaYqJrFLCXgUvI/hTm8P2Nv4hwzcCydYLH84iD1Kj4w
O611h+DzffRHEBc1U1YvmMFAO5BxwJ5XW7NE+8OYaNPgJZhqBeqExkYpIRr6PeKk5WNjOp8dDo0q
ro+//INhgINQ/SKY+PPVrLgL4lcQ3DhxpFVAfLjkM7IR4RrHFumN+8Ng7aJZir1rBdo5W0Yn0Ljb
nZpl/9SpDK8uVVl8Ij4iK+aLN4wOI/p/MhHZ84mMxBGrhJUByijYF8H46/b5jawOFQKk31aJnqvP
qsK/p5+aOd3faC5WN7d69eZmvQzYKtW+2HN55mif2QZW4JGOeId2sBZNqjyDPUojUjU8Hi74C7fi
4OmaN+JOa6PKNIbivx8LAXb3Lf/dUHKuIU4FaXeFsrX7oYokA0hInxq8btaxQPrd3OkFkOpExaW7
e0ft3uNz1XYLnY/uku32DjqI1qHl4yEk3BdNxQkCRwhse20nKLixfR/3kB+CKaWGgzk/PAfOERyG
4knr/NM6lBNaD2gB6WjSe7HAb9xxlhHCvu06R99rG73F3i5iROO1vEDdZ6/U7DcztmXItyW0LHtT
wobhc/dtnfoXxGas5+DhFhFJczsjJ7glO9vt9GDFn4T0ngN7xj4VuavJ8Thg26cHY3eCdRaoMFmy
icPkBUlB0sGDP1Ix0spWJs3Tm2BYVySnTrvjYH8zFxFn0ozzg+4/F+tumIzHDNEvKUwptYo+Cniu
4QOg/byO+Mb2BdVJNN4MybMR+XwQ3BKi974loJgTALZB4SQFG9rpdFZ0YD9L7ZaeoMjo9vSmpNXz
USZDHRU0o7NFBsRPJLVGFzpOdi9bscRUWLaVrX+IAx6QpyUME6H6+GHVDC7zuNTaSv2G7mTLlrTq
hDP8gRTTWW/lwftwSVqijQJ+xcYRbytdMFGJZY6rkp5qDhgUce7b/3/FkrhdzNC6xeDcnULIlT08
TrB830U9wxRMzHrB/V/a89UsJlKdJfVyR37DF1ZpSy+/kVnOA8/DVNJ84UVgGM4JXQJy4k9Mz5zo
4LxJi4kDJFpd0NkXjjKtQz81mTkik2Bhi7KBj+2PKLkRQ4OchPpm4mB8h+ShDvhfvKfEnplvWFzq
EVe16vUXetjh9sealdetpgPP6mcBFo3un35Hz+gCPzE1Qsw6C/u6U+ddFqT2vGWRKUC4aEuSg8v4
Q2XVk3xCP2ppb7wokmZ18KIGzZYdVR/yI/EMI37tzHl5D0B3fJFDoGqpwy914MOoSWvf/AAduQbY
9RfdSSIXA2TuxFzYbgfmkArk3WnZJnFQsHLUvAi3hhocE6geJ96hfTtpQ3W8x698TPH0dTcqMzIn
072C8eSHxiRGYoRVKUgIxCWvWM3s2yx/IWPgiV3ptCnWxKisSyAuBiIurlBZC3y4wSt0dFcTZbrB
lugarOEqG7tNSYmMB1cNXDDkems9BnaXbnZ9p8UDGDYfkCYGQMWuUjl0EW1KRubv62HSwnYwa3q8
VFjJ74EV3RHygC9FWppBRFtDa0vmdyStuNcOY0wkI5oNuJWJQ6JK1v7gvYl96NTGI8edJ8VS6CxK
tckmDDMNUOvLMvHEkChbu9353RblAnwFH+weqhVaOgnQBIwV0EfSCI596FXXq3xQt5Dy5/V8qx2n
ZTs8Be9d894I/wFPRqYkytyrqho7YMxy7R9zcO032bx8GbX+CFdzGu+tliDeEtIKTF7i8PUcyEmP
3LgevH2vBBFODBmkIK1UQH2RFiK2rVJjWX0IPRPPx1W5Op6JXlIy8W47k/RmyHZY+rBj89jcLapC
NfoneyjRvEwGYuhZnrCO3wdbfQ7yJLScyOeVqF6uJ0/QsnvUJE5XWeK9m3g0ST+oqcdD5DW60qIF
YwuJYu3OpH/f1+m3lH4LDKjdw9Xg7gmgQKmpCLFeL+vRACxkn8OpFmm1kSM3oRJOBeoOwbm4u9a0
FhN2juxB0ZKxXxyoZroLN0U7DdUbDYCT0nT8wLja/qhusxYvJSjqE5mq7nAQNso4KXwXC2KV3WrE
VmcNFqY5KIEaBjNMkCOSA2VCnL0wW/C9nSfcM3zO1A8MXwCNfW54E1hg3Vuagb68E8XtKttlvq1m
F6OZCEj1MO8R80dx64dmLzs8X2aEj5SlYXvKnA+Ri6pzZ42rs4NTh1mKZRcExRJikL7gb3OjT7Gg
JqZ8cSzkCpozQsT7cxH7scc08VvZXEHI3egpNH/D+pT1Gaq2kw8kqorjgHeQznqVpZvREdX7d1HL
Zpj1nZexBEQBInYyuCo9iDoRW4xVEe77r9LuNVuSK/o/2tEndEnuzhlg25OQXBZTgEwnJV/PzrP2
k7S3szxDwJdOkOMje0PpSOOyB+lIG2G3iVHX0gg1GbAOcDlQ14NWxmEPMDc3JbKL0/spl/QOpccM
gcb9rI39X9Kdedu+sa3E8YvQ0M+b0rMETtrOv9hAziJo8QOQhfoqExiMowpGDL4Hbyo1QtelMEHy
owvJpGvm7PaD5/hbLbpvKuaJ2S5G4ufeCCQyWz86w7saFWWO8VCejduo7eDdePgOJyY/RPPNrmdt
CWm+lYejTRijM9wI/e3/2Yi8fJzhE05atoKRkkWIOF7zUG3X+lNICoMX7cLehjQnNZFpPam/V6oP
tsTAa99QnIYPU2TiKxplU2tZmcW9TnzFxchpdLZC0Sq/ul63sQOmTcUVNx7rpKn3+AlA/fXW9cRR
h0lxUomjJME4VG+AIpyYStM5I8ok0OIspYk6FwJsQ/2ftbovxCNzQ55YNHE67vL2W4cYA7W852nU
6w/siaLnokgpwvMNx4E2bAHBAeU6qeLUhIN/taBNOAd+iPWcZ9lUleeA4om9ABLUu6iPLESwBHdP
oXMxOMbthUTUTRJKR5bkR+5IsWc3ICaqmYyhQr+ZbHscepUbjJKeik6mQwUx7YtfT6mbiZhHEiVU
jMNqOG4FYBQVXbgq9DWiFgHBJT0eqVc0upb53G23ft5S4XFGP9BMb6gC7yaV6g0y7CTsuUDtr+PH
ka9KchCt7cBLvPHTnZ5BtK2/D7CT47LH48dIzm5DizV4eOP+teEEiNAg5BiRAdiJfTjHcsi0bwMX
zP774aIqC18SrUhWJ54e5lGtWjYcnp1elY+Anf41+P6gmxdsxIoE/4Xr/VqPuVI8dZpqz2Qp9njL
+T4j44QU0J7aNtXtUtEL8pkJj0DEGFsuogbP8ZJejw9lVwtv0Dl4uxIZUo3+6DWUGAifPwp4ftqK
RvJxGNZdNd7orupoTwkuuhUJdGPS0JwzKVQ2dsVSC6p4NiYu0m2d+kWDMqshWw0S7uF0X5Rtxui8
r6CA6c3Zfh1DH4tpf5I1VzMQjwmfehxHUGX4Y9U33fo2R/tuQHNEPy4xisvG+YuF+mlQoJuFHSeE
fjHVjriEXgUYJ0wLQPdnoNk8MuJNhvS1RrzW/1XIMDnFBMJDuT56ufHx2m3FIKO4xGVjSHMOX0A0
5LcRPopX0tukZ9niQtn8AsNrjr0ar/+29wTlTZefzuzImCntoJziq+cY08vmeTyw+NvRPX7K/3Tz
BtcvqvNjMGgsYaxqG4ozJLgk+pN2yFOfqLjMVRrPJqqf1EokpjOFsWNKaVRx5vGxBMwo3YzUGf+l
sHEzZoehBmk32u4dA04HI9XnDNQOOwMZYOiFWJyW0KiF5BdknuPZARu7NjaHKobWbgV4ObztuRM+
OpHPdg6/kHxowW+H3jKTl2V0U4tBYHd/+SxuAQqEXIM3xFrT8C9LifIq9JqIAFmh/YdxElhFjAWV
3L9C3sQgFkX75J2Q4bYBOg2H+ugNU4ZGxS+Z5jO46BSoxbRisalw1/v3igKGakupxm0KFeKRYxtq
llnVfxsnfQvUWDtYYM2pSiLHJtOBO0aZNRdL20GGv8WYLj+jXscVIILOJBQiP65vhEw5iC3NEkUT
FZuqhytz2csbvOUXPwQ2UjTH8O7bIAQHOSDJAop3wp+b1dywx3T14Z3KSyLT2fW1lK8q/M7eFBAu
ZSc3eRHgnKIFhkpMURdW0kkcM7/M643yqRIMUzacWpX9sZBfFdP0eCYef9W4PoPqna48p67U/ZbE
BXoL189yt4yK1Pk1D5tvZXZawFj/avMr554Q1Kz/LNoz/Y0voWzZHniBA/2mMGy6o6N6sQrzspZk
4YutXaf1hRza+m/oiROWAvh3XdJfo3ciNzAzq6botxDzUALSpf31aNckoqLDnPQcqUeVtgeYqurH
eBsxFq5GyA8cpi8fjJMUmNPzfSeeynLUancmXr9TWGvTzhQx1zPtnQxtnzRvAf0pz4PGA6QRUCcZ
I46tb6re33fIobs+t/bsHfUQzGppdkGlyCugD3rlA55VgvDvdlCRT19wQtsVKrXwJy1dPPkpZjS/
eZqFkYHF+BBgg9wzFlJB2YWbqYjnt4wRZ3WP23kZwc0NMUuEXS/8ujQXvL5kgG0vte8mqZ6PKscL
/oaOHG95L4r4r28nXoxpYFoFx4YegItB+fA28NiWe8rURTuH4txjLwr3pnUWKVaRankuJ5BDVAxc
l7+4b5q0Sn3dBYN/jHuENQCwnQm1fbE5CQtWxpp0yy7JjdGtzhJRYINPxF5xuPRKJp+0N7ow7GEH
5Ig0PGEOZvOIeD3U2P5vILln8TDwklsI+GzFs0SEh2viLvIils+TQwEypPSMgQfcBXy45x1wV7PT
zn45v7TbvAoePoEz6HDxZWzQqSJHFcqC/TigyQzBGkg6QXKHBG2mELdg6agR2YdLDaKFLJ3kboJ7
putsh4ckV1YE1CO0Aahtzhan1HSXPLbpjtP2hYMDj8pL60IayscLvzlnnj4FhSS8ISXvP1Wnwt2Q
XpxYmIPNQfkCkA5J2lsA9odh2ERqPsU+4jTVgiYAiNNIcW2jOPh/PIli97tuyP4QVIUzjnA6DHCU
UUhkPSi5gbGGc/eSGEsyqO+g6cwi2MjGAte5YhbhQy+eIb/12MloezuuSd0ZpD0dUQx67LZTNI9x
LxAQrcKLU6OtpNIGSOBSKrMxkRSWhi5M1lBIhL214ls77buey7vGOn0Be9oyxWNZOoGKjGQaRcDW
L3ukHAbuIRE23HCfqMjOPk2tnVB5/G0S8tAD+AGA3Hx+fP7vkXoPaWAIc9LRqdU/X8AIdEN5lXAz
rCKbAq2T5yB0ql/9TalOOrq5iCoTDrb8PSuJAN06cBIN0uvycGcsgqRzzBjc8ePgjxVNX4wk4P1r
64YP2S9DNHmg0RbD9jhF3izdaa9/WuoFdmy7aBItERYnrq87m7+UYG8XGU3QR6ABjyaKrex5Wdr0
6M8WSlsBwQuw63VbhvWtl33NNKR6ymGNeZ2+mMCY39jy8N1JjGlp/NnuC7kFj7byiBTGghaWwKLA
FXSY729NNQFhiU9ZmTwzkGGCje9fOP0iv2BMFpeP7yepyaFMlWv9GlQjvB73pT2zQJ6jGCbg+JDd
LqS6YcfjmuLop6H31LOulDZpU32N7+NPWKol3io8YtqqmBvKXzqN1YXxYeisWvm+FP9NeTkUv/vg
WGQEJGLhxbswyh32eT+YljreOm9T7edOkpZud8F8lLP1O1Q8ppWAiZlbed4ADw+HJBalGEBLs2fD
V0ABzVnmUceFlpN+K8ctbHaQ2rukQ/Fx44YamBcFgugH7oxKuWpJvtzf5BI6L59Jc8bitqKPGvli
IPm2iz4kERc9fNImCjMLVSnGFvP4iZWIUnbffzp9KY2FCvyRUyU0KzKvu8xs/766JRFk0++GLOBV
RuD+WwbQ57FX7jGqsqUe1zmwoX7+zEhEnsdTpVZfZlG3B2uujsr3SL+/YdqPzB5DuUfBcsMOBvvD
kRn9EDMN2616jQuxsIzMuwB1sB79ZgYCTaOBUt6H/V4k8FLCqOZXKcrVtS4mdGw3F5LAuA6HVv//
dq8herSMjw1oiS1AZaqQNnkN7W/9TNTgvHV4orqh0tdXUXCJn9smej3GFKiMNyJzK7TtBiJdVO6A
c6WUkILvH4AlOrii7lVMnzBwe1sfFMjB+sHplXCb+6y7k/5EZ+n8by1Df61ZTvMEfG+6/RsIWPWp
U5lmS8OlH0DwJwPJ6SDSlz4kFhzG6nXp0hkVROBvpHWttA2njaAXe9Mt8WQzUGnlatQ7VconVaIc
lCULN+BAsFZzMtx8L2YkUqjT4gCCDfjDtiln2fDPAh7aQIg7vsJiRuwWwVwrddnqFZbxn0EvQb3K
CYjutn7vFaVNUItyhnYvJn8uz3/Vy2he/O+eHRpqgW85pjcsmcctZCV6rK4Q5nzI9LZPjCJDvBLw
AY8RA6cXnaG2rldH3TvZwLiw6l3aCaHVFr6Xa9OTVJle5pTXdX20OZP4M3dfxZ4Asr7KrACf4umF
hoc1JAIwNGem6zuwXt4Kzecrv3CJwH72+YDHcwBlA9X4Tz/4Lxk3nJ691N9UIecpXXqtViBch+v6
VPHiJr7/hHl1SwxtFQOrzLzX+9W21xYHuHdOJImLdu0jKicaXfurTT/tO3TUpkxfwG4rx+4NDr5D
ozWLWqU7fQi4VnAgN+gtDayjNdml8ycacDqvg64g9SJVsZbBkOiTMg8Vfp6xTn7fl5gl0J/fWEQN
+NZD5BBNwVvBzGBO50Q1yOzhR9V4vZszRDmGOMAI1C+D6yMQXnlqbdI5Xg4ly633fZiFuMuK1AmG
KXnTn78umaUpawP3ODzOFGDb4LCL09RfZzIEM3wvk3ejCjS+slKn/Lq9ROnH9d0/5BOzN1QPOBEs
RwAJJlfzggz5KFPChyYjsmYHKg7a39mo3Q3GWUfu+0VKJCZKU2qsBfJ4/StbN35iWz5W35ybw9A1
VTi/QqDeuvAwRhlmB5uUDNfe/SSq6+/5jydN1bIeYIsaCeuoOmKtDL2yVQex32n2Sm7KyLqV82ze
LdnvSyShQ5Y2+nDqCNY/g5joFBa+peW+0WMhJAddksT8gYfmeYQpLE++F0Y/x4Ke8qAYy0vqlF3Q
PRpX+lOG6Mzc758UynqfI2IoIDPd9qxkoX3u36OHUJkokUbMlfZ0g9O6e/Q6/1P6d14iP3hnOY1U
Do6x123wBoID5ZNaH3Y6B3+PKt7ED+mku5H375Zlhvh8Hl1G5WZ9qxiKf48D6C/+J0kDIe2vdrem
Ma4yAHSXKNMvtkoIJ81bIiOelzNc6woO7wp4UMMsUyLJzQ3Lfr8GPfP/9D4Ut4ARWoCXUsbt5e+5
tPXvRVQewvEHODpvV14c5W/nEs4kEW9VI37dwIgrIiuFOVQH/MY2Q/QALRrT65v5MW3gC0P7AZm7
KZ2fWWSyjLXjV1Sijlurg+Z5GFfRrqm4LaDMPI7jrIMutcrqZndTxtcNBzAghqIrbsfsGG5jAuuw
o/5Mzc1PgmkFbn9EYJMAD1PyS/C2Ff9ePIKsH+1nYDcZDMGjYwEVa8T+O2Xx8RgQhH7vJbWBa0vp
j3P+PeyHZzh4MNdhJh4MbTa9P7Z8g5SAxGoy98uz2wcSIPz2arfCAC8E5hU+pgl+/cU2IkHw3r85
JWKIPsqI6wWO/k7ZEPdqChO33jACCjqfblPFuBifcfcje5ZtWhZxW47tVN3uF0R9n1MqLI6ymWLc
TJAA3c8KxxYZb3HPPLzDH8hymZmwEeGahDJlttfT2sAAZuPR/hND6f7uPwYTDvdeCunlAX1Rz6op
B7HvClyD+Zc+h+T+2Xxc9UsdQfo8ttcyrMS8GyMftklCVTIxnaIVSwAsgQB2ptvhpTQGZmO9/mPF
VJ+xgDji7SAICONuugmsj+ajuX/5kFQP3QrGZp9V3jjmZ3LRVOntP+ZSJZYbV6LovAvIDBcXY1Zr
zSnmD290kKmg0jKPA8KqIkcOSUdkjghX8ISD4WeUQTHBag9QQl6mtLLKesmrEhCDebmyceN3j6Xz
ZsvWlAfMBGv4nNIa5nNh2qgkot2cvc1ykv9GF+CwAB9tcLn+D5GURnz04sFRUWmWTo8OTht4AvDy
zs4vwf8uC01LafqIdZg3zna/2yswHGQnwp8sGsW+ryNgVG3z/XrnqoghhKbPdFBhcMFxccn33PhQ
nG02CqOIrOyqlcgLOTsqSeXHDwR94fESFTEjeXkhXDIv4OXBvz3o0ItwyKSpuXxr68zU/cS9qiU3
B+6rI5c24YSk35UyjJxvlQfG7lxna7lnLk+lxrkBRhfD15tatI+R714+Gm4lHugktLv4vQ5Job5g
qHuDrcx1aSCYl8YNTUjW4Cc9wXS5ULfR3V24Yb0FibGEnefSdvdrNEVP4qu3JgrKA4XmA8Udhz4u
pCLuTtYRUZmlin62OTB7Jp0oMz5Lg2whHUPDAX5mGYv1qBIksa16AWTGOxkR0lcPwi4OVebHVJoz
VqRoz7QgbaaDVNLN3FUQivbq34XNUQDKU+BrpOvog2Q5Nh5/6lWP4qVDrBf64mj6Fa1PwUERXUMF
YOPvTbvdcOVWzJI+uqMUGleSBtJ8hlm493cSm6li39KfTAqmXL8c+ukDTeMjYw6nychQeVCGlFWy
LZjBifI4xa+tXBgq1C8+F9eMCYiTQGr2rPdP0v7t63G6spYbBvrhV88qV7V1hVQvezx1r+WHJUgd
ncD16753N2hl2TxsjpfPTeFF28K1RbSW/FrCB8ENCfZuYRGW7kqK2ilD92PxhobHKESOk/PuWHMX
l+QFyVlvoPIeFOyhCgk9BupRfSw6CVHjiidGLHWq98rsA/xmhc5JjP2tce/rIh0YIZBwg4/GJ6np
T0Aswf1BWreKb6uuI08cjv1NXS0NJRlSSh6cnsswtm5DbcQR38cyVr/XlZ/KQSDejnD+U4PAn/Es
ZSaQGKPUqq5PvRSsTxwYU8iE45BTM6hlpyLXBTwVMmwnDKYVpRD/Iveyj9fF3H91rQMC/P/npJhj
yrH7Mqal0RT7xqk9+wg06hqm1U78JZn1JrvCWhrp9PjB1Otnai+V6Ps9jDbiTGAq8wZsbpRYheWa
ioYj59VWN+/73jGLNqqIjh8BtM5Y2mpYMAQrUGUp+qV7CRGoUWUvlmIq4XjhuGeDEHSdhjE8YJ1n
wWFFImxjYRYhsnnNl7F3kJIzcPN/d8C94HUqRvAO37Nv4L9XfnfBiUZP7KKUoHm4Y7WDTGSBhz5w
t3OZSVz3tRnSbH57BNd5UhVqzZZhDJ6+XlDFYTQVt2o/pW048jXABSoF9ftXMZayWWU9WZxoyxHg
xIT40a/X/fznmaLN9jLAEQ61n8or9+xU6q2MioR1VCuwKHhJpYBFbXJh/Z0BrM8t/W+dqvf/hlr5
pjyTNS54mzzqRlaw9EMM5qbzruTCC0s1QVEd5iTqnIzbl2QWK4JQu8+NcVGrDuBj/AmP+i8r8/3X
uiIjDTfXNALaGDKr/mQAmpYAIkpVzVa4VQ9a0rmn3fcC+PsQJHwd+bZmUsECH8xVDg8mfGK8eyhG
wd3+2k4kCzdLzYWurO4nkfMO1T/1EgYIR1JpPTrG6fa+qFa2AYHWtdbzYXp2OQJs+n7uYBIVtOMR
0qV+T+6ODNbPclDv6pPOKtqWAoXyKsUEuFqVXk+AnT7U/iwQEUN9Quxlkhb4JZrv+v0AeAhJSRc6
GBEUStLb3kD4sYoFohjc99y1AG+WOiSVea7uSIOBZ6cdRvPht7et8KlBvC1IJVWqLDeWDbCt2Y0i
iICxLwuWZap4XMO8fZFbLsdU78EqYOAkm3DGbGG9wDLmMQb7iMn7MIfJ/TbRvzdFcJWMWi6pqJ3s
VbDSnsxQkAelgGT0P0NrRlFoI1Z3RyjEq9epda2P+KolloJ0dr7H1DJLbld8yn4/CYlYW7QzdRV7
i1X3Eho0fhfgHfWsEagDrl4qhzH+MvzBHjA7wcXpju/x1RupUPUKXsbr9iYBc1HnoSvn2WugmxaO
z/SK2aV7IrkQu9oPSsZq1YbC25gD809myAfa2dnvEc4BZcA877JMg2w17vs9WHtb9aQZdZbf03QK
piQ4Abq5flrH5SUZJoo5SDQ+jyKLQSaC4fzA9Tvju93NQGwWclPkvWCFKSpnk9p/lkgXjsAcmatp
ox/fzBTLslVSWouVRrKwX4nhpjnb9bxWkCBIrcTlOBTLsqM72TjpblYkeiyGvDqJ/S1MdtuaJBIh
A88W6b6v9F8/DlYyOMEw0Jd39eEx06xy/7UvVUk6QOjzyEwV7g06D4+uDG7hw1qrX/aAbLCvRdvG
lrVee+F31mfZhgltlFsnmygsHo0dtt1VvVvEzJrXkcrFxjXwZXwQyRuXQCsp7KderuQPrVJthC7C
WB9YhjYEsbwvPs0uK8IfWe4SL0zoVP26An25udo7KGmQ9EbLuDggfby7qWKJx5jzMA4tVFYstzPB
Vr/I2T5Cr+0QCoKVC9fSX/6OotBVPEWmKZRIIItDmrGCNTAzSBeK/DO6349UzXT0ubHezilUYGM+
mujeaSxXkgYl/cCXOH6Q7uLEgkwUZy07mqGN3cYFAlLuIUmGpu0RYnN4QdYyMnIxoG5KbIv4Phbe
ph5eehhjCxRXSJs+H26lDHvIp69ftH7qkmdmxqhwgHIMw+Z4TJL+DVRNyraTI+RFmXn8t/MbRMN9
WDEL2oam4ME928kXCA+q0HJN/WM/Jf6CKCEk9fZYOxQVmiN2f0nmXMZIBV8sXeqwbkvyG7tXU4Sv
JkJbqCSDRNsigzsBG6LUJ6HRmYke28i13HO69Uz1OJQ82E1fAMvaqg1HSLJK02aSQZhXInVuFjdG
QvI07dGYiSuCR9bXND7LR61kxHJiarRJAk5KZGKwf+Nc43GQVsDwqr0W/ZI8omIQWPdt9hkkH+ka
/9R5S5lE7/mg0jpd5yo6b1K+UpxjYNLeCKon7K+DzYdeG0n+col6+yDYnp9p77bSoLNsoIq5GRML
96FktdCHVTyNdD1xUO1X9nlzfXFR/TVU2IcGQVDigK3TV9gut1brNmUvSna3BlUkONUPKFpRC8Im
LRdOjTrkZYrlsosEmVvQfIWDvwaVMq1eCFo5Xa9nF6f8Lgi95YBdJq5UuTFPAx/77fUJmzQkYzzX
BjbUBDyH5MjixcySl8ZJjM/YN8NKE83Kw/mPx4Sr2ncX2P6g0QpGsXf3ZVR68F6jY2Xj0JSifP+p
CRgr+abjmH68wFFizCbLbt0VRqEma64TjT4xL5vlpfXSQgnCflC7+N6OvnKZEOeGiNHN6CDTm39j
p3fKHfD3AD7PFQEluNgRP4EGvWVtyKWTEh/oby08Sb5EpmboZ/PkmdYeOYROL5DsXn5boVL6jXhY
QF0Mhw4pAdgS8ErymKeB1RApXC24g7O4/W1pFzQxMVSO8QBu4jGigR8mlIXmfVxS82+6x6Imk/ix
2YkQEaETeaN+v8GssXtkK4iqPBffUzXAszU5RPxxZ8YBSS7pd4Ha2jgCWDf2lm+1pGD+lYRqZFh2
SHXki/Q19khJBpTnOPX0bPPTgdeQqWNI4TJwX7ybJUfCgRWfufiPtN0ZNleZNbxXEHiGxdyMbk83
kTO8erBOnQh0D73tPdysPVqLH/9xaByYNCvDNAesUNn7YsPlKefUyxZAX2N+hVgBuMnYc/84UQLd
xMi68s3hdGCAxcboyxZxziv5JHavLctzTlOl7pHoNtButLTnz5pC2x3HIetjJVF40PNX26RQug/t
6M31bTjwFM86EYjCMpNiLk+0y3lSD0gPD/ElyxojDB5gZUTIFdkvKbM8exUQoHU+AcaFNuWZSWtW
yhCJzC2T2phtM90QVJgn3YWfpoFDhXZ4gO6W0KZtdEi0XRxDQh34ihDrW/+DezfQAbKKxtrHQF2m
hNvX/QbBjq9OTR7Xdy8aG2DRMakBxr2dOCexFthLoapigI2bP2aWoJvC38L8+/GgZpK2R6lh91RP
FlerrgTV3GF18JAyGIiYg11nflQlke2uR7zxHgDByGA6DLLyS4xQXzPz25PHuhmjaOMN6hGL1Mgo
A19wHjATtS3PAVwxLquOCHiEVR2U+7tnZTuYeJVHxGZaxjAxE2QcP0ky/zjePc6YnGPd8Tw2oTj5
Jr5OXbIOLRrbCcd7SA18G8CPV1pcNbwDXEIXA0P9OJlDsCWQnKIs1qjqqTt21fcXcbCz3uFj9bgO
zzE0yeDHALejHLHxdBO6pTTpLkdFYsmH+5A9fmIxQ1dAnP5gV50bnXfiUlnT4c7mRCt/FH5as6nW
MmiQ30uGKt207JSb6HtMHTHFy8KKa+/BTF6uF6X4jC3nAhAfhGrQ3BjXRITRpWCbzlWL2zWh6q6T
cksjBKHYsVkPzF6/bwOn0ts82EwleCk7IdJJO1B1I+e83/DpAQakaaDAcNNxpB72tOUPhJs+RByh
7XFFTFX0LSsY9SUqTDOlmInEeZ8cCmdQ8U7M31+5ohFB5/YP6tHMKqWSIW4AhNWc39qo009zIXh1
34eO5n+UlZqF1h5IhO+cThppu/BmcWj9jV/8bHNhGT15nR+fHBRI4YWlBB0+jws+0v94wHZttgiA
IBe8jxxqx/n43Wk5v7vFJ0ze9dwg6gwwqIzTq7KwU5uqEvJ0WVdOwq7OP6FCafRcGj2iHxDSCLKA
6a7HPaip38ACmOB50FDVFrxOofAQYLBsDC6jnaoRX3gsi7clwKh4HbqMyqPet32dnkwWTO3iSIW6
K4f41vZoXQcEdgqrkO3I1e0OX8IRZhnaXg0LG2MQWTqPWlp5BLpYYEWO42iuzbK3w5YrNGcvhzSJ
1Oa6l28LOqa0lzmCz17ZwM0iZu6OYxP9TBqz70humYt09RUBBrG2kqD/piXDjvqdsNdxaQxEBq93
DUZfCI8nR2WcmJR4eOUhv4A8Vhj6QM9hsHcp2bgWwPsgpi+MN6W3z1sfdVsAimd/TsgXACdUSLG4
Q2KwcdMq6E7VyOzZkEYoV8jJqVbEFelAfNrSHmBKPDAURM0MVEjXpMG9TFhEruYhg7ShC7WdGJrv
puHw3osNeXDMv+kc5WZypzDXgN9Urwg7OKClvlFH9UA7warElPLZgpm0K/hWbQBIEkMXzttok4vV
Wj2rQxZyJq+iSBX0k8hd+5JXFGOwl8N+1rYyeyFLJEyUH4dleIBoXTBtVSVWFq68YxVmMejVjHOv
fSAjpKAKBL5IxhGzzKYoP9fUlewCaADrkx7A0d/VOxeR5FPqMix+kC4N1OwOFGM1bfgMKSvPj3Ow
O23oByb0CQiynWJ/divAHo80loZeM7Tq+iHBXK168VWFbQFKchgFsB6P5KScBg44Q7xgnnzShUQT
ODs7Z6deZ1j4vOWWuzRKoF2XKuq3AW4FPvReCify74hvRZY6Ap0DCvb9kfEVPAT4W8/7SEHVJdt1
ukk2hLkohWtMP8NevnA2NIH/Vd3sVAe+2mtyXTwD8mEVfHpfYytB99krvEC7ZbiUleGtBrZcpByW
j9CBm8NdXNE/lCmI32JfwPYbdTmdloMSjyC7lPm6uMdav58NV9FVKVU113i0fqOUEPU1n2pvyKsR
Hj7aNOe9NTY4VAVLxHsMHwZ6lLtnWQvxhtcKFXNzaZOQdKiGIVpLL9B8Nf260VK1HXCvY4r260Kr
W7CGXMiHsP3JH60eC/cM/jpSa8PsMc98+6GVnfNEz0pSoXHmiU3dU/mFAh6WmI/vh7HZCg0tJ3vC
sY87t+bkrkJjICE0Njhf+3C60bsGiC492x/jJHbnTLAhyy+c2IABc0EsW5FRg1kiWTXGG/LGJBCv
BwzCcFXdogwoS8axYn9c5KNd5++9vJa1JfSjMG/5rb/sArb7EGKXqwoT5ui8cUn/zBFCKZiiEo5C
1b7DNwby1aqnUYoODqrux7ESLXBio0KTCWIBcXeOcV/PSKl6uzGtTe9azvsLtq5pvFkJeeAkx3//
bOmvaktWKW3ZimbBXmVkNCYGEBA8RlIGAwGo68Y8tD5IRC65dXhY03aZG/fy89OZuVaIvRbENhVu
45NwbNNi7eKgQtfNNJ7rN69IymLXEt3qJR0Kmm7Nc51OfJcflyAbeUB1RCaIUvKT6BH8YumcEviQ
Mx2dy2xjayMdYv/EJWHNzLY9FbHBC4chU5cFtr/TaUt0M1+wO1W4TPifJ3gg8/0ULdikAQhnaJMU
sA3S+08Q9EdPR9yBD51FW7cn+sv6dQ88ViC3h/OEE8o+yS9IMB/Q8cDkL+4bY+5ocCFlGOWEpMdr
2Ra5n/6mG5+1pfA5rCS7xN0FhXcb9LPcQ5/3ISbshps19fvSmrl8AFrkvTGbi1MfPACLaDcJz3ur
HJ0mq4BqM/VJnA12+FspGDTKx6zavh45hGKF9QzJnWQekUiq/qEDvYF2ivjiEceV2PrT0aUalLUV
skZHtar48hGmObp0N32hhG+hQn/py07klfLXhq7EPqRJ7ejIbdRS6ihdSG5S2LnYAqXHXK4WEwgd
T2dz6/tmxezIpBA9fvOAUQDrCacS+g8Li1rspAI/56TL3yZiJVDnnr+pdD+qdgthvcqmgMJ9M1Tv
E5yrfDNRh8gcZaavcg10TDWocFRE5FtL7PGhXGiamCQbq817Un0LlXHNcoG/GGp/ZJ+/WZ+EmNyp
j5m9jPzXFYYJMFJ6NPj035ZjO60iAWLk+/v97YY0V6NpZ3prhAG8Y76Zmsa5Mxkybl05JznFZCLv
6fuVjocTrryWybOoxy1n10PlAsJqVVhVaVZUpZ14GCZXKYjUR7XPJ/b8UfWWadbaZItyPTbLhuaO
AnU8BdTN8Yf6b9VJMhPpUs3xayaz5uVU9Jwiw0BxPWrpn1Bw3xBI4R1nekPIHvUIEPpShcVNLyjf
bNZCllhhG1xSTI108nNXVdQXBcbxcygCiyNTC2GQAdvPZXM7ah+/uPI8SlqiCjiP36xVP/xXXssg
yvi4qILj6nWFWe34fkthCjdw+uMv/fp1RVa0dDeO0bEwnRQNekbTUVcZ42K0wbtBHFT6LBfwvmfb
Z4c9tdu3enghO9Rmar77tGiqQu2gQcT0Dex+6/evqIn2deUZqFemkhCfEOObs+gVHoqjbutKBWVc
sq/xUkoQ2nqKZFb3sRE5GSA05cINA5TY2ovK5aMSEbXETlqzNBKm5Fxvi1f/cbRMDbyvTFopD19Q
ehxKx3oFV2zzMM/ltYII1rcV1wSSTpuYI4CESVECsfOMOhipw1GWX5kqcQ3qKms5MRBZfxEeR3zr
soPv8JCCcDPVBEmvaYu2nCgWIShR2HXyxshdK1rFmYCUFIDA7/aYiptbU+G2YamC/D6cVUgMD3h9
gS7U2mLrPlyJZLbyO42dfwnMqdw6+K3gtsZRVnAW8W06dloAIlkFq6Vh4gpzBddLetbEDoFe9tB/
yi4m8rsdwQJZgnsz2fmQ5hhroRl4LNEbsc70BdGkwwCGerMW5KuCfzZ8WrKJcdQH6DhKTaTr4GBY
B81UKx6L7ec715qFliKixLCB9mBCSAB7I8Fh1V1kr0Vr5zOqtXJ0Ia0I7mvI81TWXHGMp4HWe4P8
LazbAWJlGVVjEb9+KEVl6Aosz/6Y/j/hI+EaZBkOUgiD7+ny6AgrngbMTtUjThJq4Zx3H6Ild+a8
3z6tsdtbjIOTCv1jOk8rV8iJSe2kg5B/XD0VDJzsaLtMMp6HiSbfsl+CDtGWbp2UtsGT4/MiTKhQ
N7vxPyBfgaKvTEi1O/phOssWYd3suf8YCLxFGWH6ViFpHL1AvBbbb25vPynFDJbSahSOvwWV0R41
GRw17lw6FFwukCLI5/hGEwvStu9NYgRqK26MRMVRNEBMI+1InlhAh1I0qYNAC5fPahrH/BM0Ravs
QPjX9O7jYv1ts3ibpjGdCFzv6F2N1tbsOIvXLJlHsNexTanRPOsst1u7c/TeKoqRJj1FOZ2yxpgF
lBQBu9MEagmdExbClUypOwS7aTThNs+Ca8RqEuBhxwSuS4dHD2KS1DXgCfA5u9BjRz5KWyTyBt+O
Q6gMeq1K2W2t1sRDYt74up+x9w3EWZd9dM3Fz/eVwY+oBFZoKrFobcO/Rcr/Qbty14zgxgiYMeth
SKPy9q6EOIbLCeadauoAtflOTormLHNZVNVdlQfId+jCnPrp3NhbiDTlTTQmJ9OSRi7ul0J0QCnu
nXZGfxmWcrRpIOueXt/Fcpvc+j5C983gxTBf1KjoyiJ7KJiKjxwoGof6LI1V/epXXmfAsSdJ2tCt
tFUcuqvvJ4PScCGORfvRJZnQxMeJSSG6idEAwCazGDmQ5EGb6mj+30oPMC536aUjOREC9ggENpqZ
Q2xkv8kZXi1JpmuBoC4iiSd8R68H22P9ln5jcUj7bSumys7qSvjO1ZwkTRAX7jjr12fbenxA+Tv4
Oz7IAQ55mLH/GLMESi63bAuY03S59PTzStrdxxlCPGcUEkcN5qOStFbVHPTvJ/O9mKezRZ9RwmXr
gXgS70Lskb8w1U1oXFAC2oII3I7ynxO4RebpSbHFstJt/H3NlYawnZKXeMziugr/evyBJzz+SknP
WYITL+gT3XLh1NQFy2vfTg7SBljrP7sI9t5xS4jDccYzT8/ZaPOuMQdkReVS5Md7SCql1Crl5riu
0K7J+/yiFpJt4jh5XbqDDM5Tl4OqyabD7hlAefk1BKePDSGFcvosLM135tuF1gGxSkV6czius4fi
DaUl9AyhbNog7dxvW154pPTnOMDLCHTdlco0XJIPaDB7lofP4Szw9VAYU2nfaQEpaEEBBsRGdXLH
XauFsJHMa1SBNIftQ/cuTvmJa9dm0kUdZW0u0/doG9yEMwYQYieQVnDCmIurt4EE9wVSzm/7ZM0y
xulTPA0RP45cfM8SLVct7XkK5dNLD1NtJOUsyp8lmtclBf1KloG0uCdRwt9OoReZVwI4VyTMWLVk
wmPKRcqAll6FhNp6R+mGACU7GUbVqjKK3yFHiQ+i0mTTGnBCzkeVGsIT6a19OwjaClB/WOXqyh2b
+r0CueK+jA+KGfS8npbHqXke+TCaHD7syJ4+ap7zs/cuLhU8sIwwJvm6gEiq7BWzANdAhu8mgkCt
uvWcyQGIg/4gZuRQPjQSrJZQvVBaCbnNbrb65C9qtKQACwwHO0aRdoMisa9qwE//YyWxfTm+N4z6
U5aSqVdFIvy8GwpLFKqyKG3czwfscDWqla1yjdFUGzx3jB2httl6L68+L6cNGJt9wP3UsC8/Y7g5
r2xuJqdLSAAUf63Dd5NjCO37rPZb3p/rRMkdqOBVciEKLT0epggxVUb20O958kc0qGb9OtbIAs2K
4owxhUxA1D7OPPo69NHXtK60gNAY6V/kaxKp3PhWqlSYKyruqWI6C7yM1Y5RbsoWDl8r9e9/df+n
BC64ZtbMUiNtLeNJ2EyCzAIKKtoHi2voCvsTPWXXcLZPc7qOVz+Ji6st4a3n8YkBxGVXOoT8Jo72
2ldh0usJAHIiXx/FmRfkxhf/uAqO40qoUxQvj7a+j33d+7T60uITb97m8+8DMdfBWqNh48oFlEdq
GYf7rCPdNwv04/utXnEQPl07FiFZCxLt0X2IBbs5lNBo936ZAfp09GR5BkLlyA2rHOXXY+MnED3X
uom7KNr1Y9qgu9JZS56SqGB289+TqaX9GA9v+tqNxNtKeBmPQ0Am5+Rx2kFdWa+UcQTl/exMiHtG
oOJcjOO+BCA4gNhQx+/NHPfDE1OGkRMwfvflsIkKW/mnQJhSZQQ35BetIIteJzKSjTqDJfM5w68M
NDCg3BL8lVK7b4KGJzyWrQvrSpi0kKeFFDhRrLnr/JbmsQWdl5X1u9vE19plhF6j1LBp8y/un2M2
P9boUgRl+3rpxLkE1bC28Y+LsbGknmveSwA2LvmyjCpw4t7Ai2vZTCFnmzd7+7G3Qxj3+ma7nGOP
yzRRO5gHwRBhh9R87qa/qshaHV36MZHXjYYTRfaMdL3KAk++I7cC/aGhKg8aXxavKYwYVMkUueVH
J8aVMscNdRHhzzXxBtLZW9M9XPlQx0Cvgi1ndRr9wyFULUz12EBUokcNqUeoTcSbz7iiUrBPNPEP
XIoKat9/qKfMomAKo547tR6GgMFZBbCao7pAHsC0Bq2OkW6S/r4/XvEPJZIXowqlbPKa5HcQyyxu
+pB4taPEiRU5dZLXnbKzpeYpLoNfkmz8NPKypFOm77l/+drcGg5Qf0ZMDw2OLiBUKsC2GdVDTcUy
ww+n4lNiX5iFq9PpBX3So7sDbFg/4B045CsfKjrr/OKbhiehsslJVT3E264oBY/EiJ5e1Y2VSy6/
DAr48EhlImEUHQahzItDNMgR/hGRPkB+y7jlJGthvGesXaGHIQTBaH1eZa2tkV169ggBfn9hg22R
WrbD/XHn9huIfXECe6NZ0FPtb2PR08j81Sy6Xko29SjottOHz+sz+JDHWiaHx82mwm7tcxtqYSNf
4jvKa/4QXlDF0PII2yVDtUbC32W0TDptqqa9GiXdODVuAX8xVOnm2LkD4iZMen0OetUdohBCBOe4
roF9wGCFHp6t9k2dwGF5Fi2wx1u2BImciaWaWIekluuc5KkCcmBoFbJqHRcqjuW0W7iLXnCkowCz
kPrWy7Wio85oxS05EGII1vylWvNDF/awu9yvsbGid2/Ock7nPBTeW3ZVmPMV3Koi/48FnFvEq6NH
y1GRZdN4Ux64dwU3yETZbdHxpTUri9/EAnqFgntLyxiociQKXsoy7kadFiozc+CTHogeyTKrSNSu
OXoWoEQ6Zi4M0Xlr1oTMsglB5lcIFwH73HwVH8ig6DSGC2+VQCUgJk6vAiaslHPdJVPzfXzh2qwh
GQ1nswiTIdw+Y5LN/pXDDC5vEuF9qQrtqQvFyHpNsa8jXCAnxSzrWmowoVoadTpZVKLH5IeMp/9V
FuRNBEXSuzgRKgODW8AlxdJ+bPUfwawbpyd4NE+y+B5fIIwrPvID7Dv1GQamjA2PeAMaOxYG8Jak
HQT/oVrfFz3mDJMRl7j5J20J91tvXD695PHQ/uEj8anmAugxB/uL01U/NaSLNTaI18m03ZU8NaIG
v5M5QqBFB5JHwMigwW5QV/t41S3qerKcXzwCPMlq97gTr7aUkCIrlOkf+N0GK+KqM+hFuqgj6vD2
csap2CLHqWdEV8NUlSvdEYUf+2yDAOHH4bY4UjHaiwuPtXfe2T3NSLelRJx7IbBBPUObPQJo7lAL
9y57OhelNj125v08ETSmkNizSIQe3h/fF/MG20qlUBQOuxXJ1s3ZVcVEYJT3uK4fcRdrqb2DjhPX
rtDc1jAg0xXiojQCsGXXr3M4+RJ8APeaTB4B3sEdADoP9Mj+d0qSoN8NxO2bveNsqg6kh68B+/Yk
r1vZO1RUJGVx8bguCcAJj3AInfTCDz2oONMzNU56+wfUam3/2vZ+MZKRTajd0+hbYCWcTIvJrXJG
RPxzwzEFfgWk9KwLMUM8sTjN47jBID4RPqhggq2Sjz4/9jtKlgnA+wzwV/b4ZVOuCpWhCd0uE2U4
qLfGgUV24GhxX4fBnIyPqJwfVcB/tNZ0+oG1IY2qtX69IAT1C5OYAINeW1DsGWJjzTPmDVZansO2
HdWBQmPmQAdO5d/7PXrigwUq7BXN5sg06psxN6FBlC8rOSBtWVeUH7CEbayHA/eOKbnwt1Rx6GmL
z94+SSdL+QQcmKCW7ZjIrVHKqZNwTK38EVfsDeiLYi9BjWyRRSLkxAelVRt+PbjcV7WIxK7vShQc
pPc0Q36jSw0hEQ9eZA9LoVRbns8cJWQCyjqRcv7vMaBDC9mS+hms104WczPJ+vmtzQUPrrwcSaOB
JVLM515V1TF1LlTtvL8PJt84mTjyl2lzt2T32NhL4X1XSKsDHM77GMZ956NVVTI6I4M1bIygfJ4c
2TRULcg0S/QMZuyLb6nfZrHrM25FRSZyS0kUnDRJx7jnE52lNEfG8Wcc9+ir97dkMQFHKQPzIJLW
U/2eGtzUWwPkbEJOrE8Tq1N1pMod/gDp7bG5FKVrjFkvsOF+1HRoGbT3JO6D1zeR3rq7uCZifWIs
KEJTf5joB/SarDjA2Lb5YB4fsWc7pro6KhVV4750+IDov0KhbxZDzptm/FzK5L3L+w3fEEpgO0Aj
pRYk8kLNrnvGtiHYYMRhrWB7gPb6Mn5U9UQesVJmIYBEkNu1tM9s9QhuoYdQaxblhW5VJXJ3WksR
YMtEysKZz4UMA6QyGlx81duV95QJMjLmK2EYkcZeyoBVqWQa8+R6NdytEi2S9KRuU3dzD2jTYBTB
ZkhX22cnxQN+TjQ3Eue7A7tO+RzX6U4asYIwyuClwOWjlcfGFucQQdROoQwJIP7m0FI5aMk4GJ/X
E4nJhYxB4OjVBhFBbUH8sI/t2udOikgxPVsfA5NfSymF9FGTT4CQOj76uvP8jso7NKS+O5L0ok2n
o73eKoggog+9stk5+Y7c3pcHKs+U3iuuEsGrB7cDtr8MeIliQtUQEOvtmxJyNtbmLBtEpggNn0UW
WqsoYm9GXIpW5a4X6xDn96zJi0mS/d76TRYTCnz7KZwCS8+an6ybhBvNS4cE6sXZGbSaHGSdD283
7mSM84C3grdtjZAbTIg1c7OCJOYCX3dT9y+4i3kmW1arc1Do3RGFbedaFgB8vQagZuS1xrtXmQLz
1O+GWEtahR0A9Z7ZkuweqIJDMc2GPCMGgJKqB4o62UUCwvCY4IwN5QMGBL9Xj8sProDacaT3t4Rr
SgycM9WmYtWjCK7JoicVkY9siarbejuIM2Cx02BLx5l+kPyuenUBR7NqpvdLlCEYdLvVPdDaYmCx
peqgTGEaTNzAvdSfDRGOmCqxjbnyAitbemy8PqqfLhA4YtAYbeWSdUIuNz/fZYLsgY1nELKpFBY+
1DTKYyaiXB8nYx63w3YVS5scA/+yx0yWauZMJPiztKNEgVtjvi/+2iayh33ssS2f8SR5LM2lGscF
CYMJQIQo/QkmVnOnUOHmD57moiYx9ZBuAywjxnLmkijpiuyVPYEsWmhUlBXXpG1ayGLXlG/W2Yme
XdEQGwz1PJVtMMkS4QlSADyX6yYnADjlZt/sooCqLzghmXA+jjyS3Veg71Gh6E7Hj2+F7JPSI6Jl
EvJsN1nhxeXejo1oBkoSh/tJOk0kcg67lcC1+/m/Z8ob2OWTU80Ocl0X4hq+YtH3MtNMyxGAggyk
Kt/iGiG2Ew83MmoZkxDyOOZ0G5Y/uMaU09m/zH8j5Bu8+HHMLMj/csfT+bfarYc9iHHRdv2L8cxa
eocFsluv3CBRGISkregzqhl1pZghnknDDEep2P9qmfYzjB905ZSE8Os4Sbe8pXqUJ+z/smqMXWOv
z6CYxUI/9dakLIflWBWfvpASZPe0NJepOngNeCYX3wVMWBC17Ty06auJr3OIEBIxs5WiyxFS1VTe
HEcvfmNPipH51rO8ILmgTf1xGyA6YKeZN8GwmbUYjb0ybOjov2ERjBZjh3er3ARuswwlX8SpUcA4
/RfzEelg3WaIovP1wxFtON0Z2p498SpJpg3YtWlM6QWzS60v1zjJIQfv7tGx0lMCdREc6UCSwsN7
EjSA51Mwt2jMKub5cGA85JN9MmIowyWDFWe6T/DRI9/4Cw5B1pSgAF2T1C6weg0qKZrv2zlE08IQ
BwrLtdUpXpGyixDCQ8szHx/QcAyqn8RvDMUTxqDvxJdY6KFEoJfnK2P9wyJaGtml1er1eD85/4uO
22laibXG6ILwRMEl0hCvnF4UfRWbbOnDRuYfaGA7H90YF2ZT6sFQdMaSpHIUhEzEAI5iweZioTlL
LgbiaCEAz9A9bzg4Un2wm3Hmd9vyNLps8f4iynoHSVIpzBXetwwus7X+3udCT7S9OIpFJAMYngGR
ARnEpxLToUpdyljDuBtgzy2J1OMdkSIGmM96+XcQcYE293X3zFGim50mAdvbQf+qdjU8trO6lA+8
2zVNCcn9u9e1Z1ji78Z3T457JSVN4ceriL10+teKP89iTAr82YTnHgPoP7ZRAXeRZfBdhIPr/WxE
QzQ4jVQrAvRvIdmiEiX9mooTSrZbsY8SAViqwJx02bA9KRULipY5EHrYyBXB6swvHq0Awh36MqJ6
ArDK+aCYvMOl5gxFGAQyjLCERDeKwnpp4lUxJDZ4Y7cHuJeMpO/HdUEgUdGg4urFjglO/kHlynUL
wfSmrGcmOBY06dB8UhWMJWsJzrvaMVMm3AjMgkbhgTyqGrZrfkXpfuvC7m4vrGOvNDICV0cpJTgV
weGzZdUwSyktm7bQef/dPKfErVwQ8gPYwx2Swr5U1XdcuzktUC7PvCWDKMo0tec7/JX0LB3XJ9Dx
jl3vhXt478Km6IcPgrJxa6ZjnPS8AkeU91wIZ9EqVGIY/uvfOETT3+sStMJ4qP34llo3dUKjMNLO
WcFjOiwEm/VyggS8I62LRKm9TRnzxcaO/CqZb44yIOG1cQFQB3s/9GXeMY2nGZu01iIypO/qc782
Eqv1eOEGLB7iU6uouW1Kuz6vUKHxzQugnCvqCUrMn0u6oeXaZwFkkxLvuWZ7U/5xoCyoNfSGdC6M
4z71+g77csLlcn3sASeOTVUgw5jwPSNEYwZ7GZI/uuT3Zy/bwijwbodfcUyujVHNRCIkUNMlIJAI
ClY/mjvbfGvv9psebrygvTapLtASYDWuKAHwDDjQSW3zYxos0Izjtwel/u5SYwFuogltxNl9JGqD
jUOryQwcHkNq/1r4EGWj7ypAblqk8B+kf5j/fiDlpmHrln31ELPNsZlkCznh/LWhHP26RpwON4SA
7+h5lUU7ikZAXl1oK1ad2Y+AoLKv2lu70XuqZRM1e6MwWABYKI1yr3nHcBF2nIbrZK2AQpIejIC3
zjOvQEoa8msg4vbLbH8Ume/28XGmn3sV8hVdeMOe7XVRlVg4nJTaskxipvoiBVApc8EtkTQtbuS9
BEBg8cQhojk6tCXOMMLXPctM5r1zeRW+Miiz+SHAXxni+9PDHQMOhPJP38zXvsNtx4YgQTbiDV5Q
BiZiBm2bnOGrwHPL62oYYmPUK8t1QoB69PMz7jx1O12YUhbCU4bhN9XSBx1qmTaZ10AfXj6q89e/
ZHKIdV5ykF2lRk9pH8rbKNNVB4y1UhhqKvMTINrjc8KkMnjqTF5HvJWgr+2VCRiy9C4SbcOEbBil
7I2pVnhn7VUOTW3urY6eOzw+HjzapCfYFIAzpvPqtH7HERRuYMzN3NCxs0PCfPo+jdwwPebBnflo
0uOZPPVzdXRWN2qmJK+euofpLHxClLs6xss7Tbvg/Ggyjyb5frRBjF65YVW6NIGT0+6W5NnUySKn
V5afFKDtmgzItSXhy17Gen72z2okmykY51veyAxFpijL6yfLTGZ7cp5grELD8xrKT1yogXjmlsGK
SLwDgomytsF9WF/c7wo07nqXDSom2YQn/lPCntjijKLkLE0oxze1FGh6bMN0IkfXwYEtZ2ptU65E
oB+OYlcZRBMmhOSaWEDt5SRe+Dv2hl70e1D9RXcMvaIdQHw6g0Y/YYp87g32sFRz56MhC/tL9vSl
IgLNeb0jss2FJoZzD1TsILpjHy2l7CQ9x3tIOkPJYN3hMrxDrRi4+CMPnFVUH0sSjIJOnJrfQkrk
VavEXSABlg3qb2F+LWBPP4sPn0IphSFLyuewt3QeAwVnxpZ5YaV5OltO3QAwz843XG9BoACwzMUZ
NPmoFH3JzNudZgeASbWK6Gl0vgnmQ9xr4/Eo9Z/c8XnD7J45cpSfHKf+ya4aYLRU377Zxu8XBPz1
GYbeb3NIUpN7+T6Bw1oLUX/q/VhikDrCWT2+rAGM2btzuLhJbNM+396KZ79cjXelVe68fV619bjV
KHo35LRFHOlmKxEj22Makl9fJ4LSjj/qZkY1cyWSceA+gK4vdG/MlU+2XxlrHt3CaNj2hIOufdD0
rAZ1OOt9IrsFPcU8Qf9djVVCceaAgGxHQ+HDXm8oGIm0nxuYQG48w4G4TxZNwVNM0X3tO5gQK1NB
LG1f+YkO4IEPc6ZP3rKCN3mtip4KdFxVhlLY8czH4sd/0i0SCdD1NCG+tJmGQHlN4jHeYIFC+Miw
td0xy7Fn32GaRHKvaEYKv3SnY/pFGnpJpBSvvYkBgtcm4vDh5WPuY/cSuT6f1jqtytyxJPkDQR/F
5/OpkLTYlAs5QHxTt7Xvd0HsU+PdVqJ6ZBfooow5psOu5Ekv6kmnntC8ZessM3gGv3iKw7i/v67K
E7HtvkePvrNu535DMVTLuCG25lTU7VmsSTgp6t3lNkg8JbFxVIPuSqY4lStSb6YIS2njoZZ7O42Z
xhw6pm+lbx2jQoNQ7fGpBffFJZD7OuD7XnWOGe6HWvK8jvqlzfSp8ahGdxzdP5bDIDODj+V880lS
GyfHkWtzmqgETu0zC6rFCBHWETEK+4X0ibH33VFoyur+J/m9R59Ntn59X8tDMrDYbp1vjrmEJsYi
xdhAZeMue+8rW2NTsxL4+L0UCn5/l7ALm0OMTAZth+ySyYZFvCF1Yt9H7s3GNvhmXbkKNVFmDYaF
9wh5SK5qMv+AxXoRoJueN7bB7WAEc9u3EANCtf6tGiy7YP2OT+nL5fLqp0E6qW2nQXcyGyMNIjtC
4zPCouPU65fXzRsAGeW/gc72b9sxcQao7Q==
`protect end_protected
