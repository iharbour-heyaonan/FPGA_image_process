`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
PkyhyBb59EPgq8kANKUgNUvJSxwVgcYTKLlfXroHeM6zPnPHm+ATuJPY2OmCojZnDY2A6SHiMUmx
ylnsx6jVAA==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XgKClVpS+h3z22aTgNZepCZW5Yffl4m6nNLRjY88G0b6Og6dF7wA3of30X3Vr2BKX5GVSe+jeu6a
q3D7Qa0T3sEnO1qnWdbom/P31G6nS7/pQCPaLh+suxznQX2imRfhfTkmY1B9wExxZtZBbss2GPfs
EFGX8a+efiUiZLAKaSE=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LYMHL9qwz9VPPAbHAyLFK1YM6t0YBJUbhdak6y3IQta7KscLfLakFo9QXv7rXKj3R5WEjx6Vg+9K
QUgoa/uCYy+n2t004DDpVeDamNuGIrJU3WXV9mo6tEi21Rm+kIG+CFgVuqLY9JSjwI3dhmEqYYtS
wC2GIO6hKaV0keq1ldvsRFBu71kLY+jczboTe6EddpUktWp3UM/RqnrSfHPMlZWhHp1k3YC0SDq9
gvcPn9DB3vIjXgn+xRbyzZOt/j+s8RfjF446i2RalkF5p/den9o/OMG5jmv4rZKHj9S1V3Z2UuL1
c2fxe26sNIvZ7tpz8RHVWRMloPfcPVakam2zhg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BACIRg239ZSAZHpsLobWk7IZyWSAM1rsaZq5LesIgnba07iijhvT5s8WIOIIgHZs1XEDKelSnU1J
+5cyEbU9WgPZsja6FQEw6J0GuN3L/1QyrvmNIJKsNXINx7R+xaY/n0uby2eFsFE9luplvdOyrCEw
eK82BghXwPdasTT1ZUgKiycyGYtNsp5ZaPIWXI9ezN9oHowcWp7Mn6v2jrdDl4lzJuoHgqRtkZvG
7GqevJFheGfXkRPuQGkNK2Pk6XN9woSB1a9C+FUsQBM5MlIE7zrBQAjONIQj/nd82Hlp1H4PRxBW
1mmFP7PskMeNR2hH5xwkvg4Q3IfYBlw8gdzneg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
vUWbACu3JL9XeVH21XChN1bLnACIM0U/dLRQNf2LGaDFNW9CL0o3SY9pOtV226o71+9Eal6i7P4l
ht62RU2AHTweJsgWkXtQBI0/jHIw4/gxbBebNbqZM6m3qjEE5blPsuzJ1njoX2JWCJElO3p9FfRu
uHpC+4hYoccdFayGku3vk1gwz9lLJ4FcYG9mi1vLIY+tzs0o83THQ8dLrg50Rr/r2n0Xf4hxWe4U
tJ6iUOYBQUYjeOwNQOOxfjv5PKfLIgGA2WC8sJb2GFe9MkTDoMAo40nBLK0Y8+klDIJTyx079Bx0
wdRg2JxUF3+TGlXW98+2/iWy94H1CPEVRm18FQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VX8rVAT0l4oniSvb1X0sblwaqcWh2XE0oCAZbC0SVv8fCy8dLmmtqBzFq3w2V/7nyMmJzWKNP/yV
0GW7ICEfrGaBejU3VpwaHA69xE56Y/8NSHGlZOhr390/5/UqELcFOknZEPJXMLpeKjUn2ijACn/u
O0myDIvGFiUyRGWWYKM=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dlKAt52rb1rebbUvCxUw/pmWR03F+be3vApC1VuekYTvk7BFt7xopdHrqsvoU8rgaCBc2wuCudx5
nUcu7bKEyHKFc6bcbp6J84c2uG0ZckyqBn/OHRMbmq4Vbar8C3ERI2YmcbL0Q0fBLzMosVarF9eM
+c6VfE9hA5lx9qpwFJhgk5v/yx6kjgu+kEnG+xsdWrpKrj8LIxxh6gkrPOn+jQtKQSX3o7q35Rcv
W3vWLRYdH+pHsfJqCdT0wL4oBTLa7ozdsufX9l6UDgT4ECxLf7R1TtNj7XA1jaaefThL0F1AUCjF
5WuhMqBOotpDZUmvB91yVtbXLMm0r85tK9b/iA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26688)
`protect data_block
POnT8UXZ0In/jgQnN7tvt/KAkb4n77xHpqVZ/G2B5ycr4yJFjf8rniQ4/eWDIoerKqxPkPPkjIds
bfgVMWZObEGsgODGzrTmlkuaZvJxTT0stupIODf0ZQUtMhQXcFy8lO0fdHvvPnXH/r2scUNfigPI
vrq/TOmUaYww3Vc5PnE7UAsC8zZ1oUjaugyY2b7+hDloxtmEkcxbYWpf7Ku7MqVn+VEvHULqolQt
JTQu9zDO9M7+6rGoqqw3wfSW7ireieDd402d/fEol6dJ+/5fOsW5Xo3AGayEPKwOA0BvUO2qH/4W
eERojlnyuZKIKQpdqwzLBoT0eVvJIkS3hPK7bBJ/sWu4Qsl/Bu9A0asup8scxX6CaxrEXEVXwfW6
ZKM1kJ/djdEBxJD749YoXb/G/5FjG22+WU8xL2HqqY7tFqbqoUjIRcEGYL5lhqbYAWL3W+zQNnXR
4aXQVXCSfnIqm8Nw3QjnHyYwnRrOdNSN2wN/g9CwlpRFfZPhsVdM/7MYmaJUeRAo7p32V016eU47
/xBZ5OSO0XopULb2QNd5lg1daL5hZ+mhqAYUmeEtZ5canGku2HsHVrvDtefZap5HHcxRgDq9hyEh
frS+eK5B1leqlH1W06GEjiQVeHiSfeJiHrzmp7qqkMrPzTAU/m3hOjsIRfaXwqzj/Iqyq9rcVOrl
pWTccP//l81OucFCia0IoL1Lf9BBNs8Kg8I6MOdUA5XMvE9S2mDL1nY15YnjH9vDhHcC9N2QAqux
a5V0fL3O5x6gQaCdhbGHzc/hhex6hnNVKDjhJExGtbUP4FV6AIsDrm0riVmg7DeOrprbVbqBnc4B
kX1rliPnVtSkYcfMILYwGeO+gOaGuAFQF0ZrmGgaWvTXwAHpdkyAcvoHLXrBkuxZuc4ZeuJiaABs
pW898SrxsL/GS2WKjN9ktJ7yU3kPjncUOd4iYD6FnbqHSYCU6lWvnarw/QeSuogLhf3fmMh9WsMd
Zlp7Jd8NOIV38oSURiY4qF01B8nBt8Sb54igD72kxgv64IRxAnO4j7Xkn+Je8ecTSgD4B81dj0wb
rElx5uEx+ghSSg4vDDejqhWFq/6USfpZtVJgQ/VvBZHwE8YRYUbz9WhSxnoIA+AgoUXemLtcdmo4
jYzYVEf5j76UB12YrnZ7YozAxcJ6lvz0q0tJdPnwJMDC7G0fEBXr5C96MhaAb6BNugpV1qwPt+kA
JzXPqqTpBrfnk59vHvy4Dw5G+EZEgEsm0XpjZfhiAQ/c8/BMClOJatlii/Fly7sQk8ojA2a2T78C
HjixzZwNqAzIYUA95l9xiFtVf0xZK46iy+8nV4NtGQGi6tguDuRj5cf82BiKEnd1e9FDQRBifRbM
KITTtTyogFn14so9qjf5f9vF4m06Qb1/V2NF96+cMv9H6e27Hob6dJ9S7sWK9BJ0sOwckpGjM/C4
BVGj84J0mC7TzTaXtl8in5V7i6hvM+sdcmrDm+OdJDZktxwGxlDh2mPRw+I14hpH1c9PBCwdU1TL
mwqo5nLvSKHygzdZi9PTpKO3fchUzbw0F7cPczqjOJ0lJIJhOG3jxB2tIUSJKez/LlguiqWl6r1a
aRdfsHk22gqfOliaO0lssHZOGFzlzZnwxpNCxWNtKo96FvZyTxr3xRWSlAkCeC+sT2E8BvEOTQah
2Iu1MQMljVMS2vSn8XKZnYM79p9BbrC7vHO3RkfKKWCH275EEXdK2MAEakMZsa8hh7LVyTnWCjcC
0LGIE6K1ArXg1b/hebZc+q1PcpZBSCLzE+gfpG/QYDdmnz0b1njboAd59bafS3OFy7Lyr54TOpdg
Bsji6UQDp9hMlBT5CU8C61B77cN18522vv40hh6JCVnG8gtTucOWUDVoNy/7P1gvj+9GokBwwTL7
tASlt39+2mcHVrlz5Q3Dh4bUKFoG3QjYXJhFLxnsot+AiX5kgAdkO/E//apCtQGie45ryCIrIf/1
elMiZmk4cdm0jXe5VKxh7BFEZAdrM7OL6lItmjhMJ5IfgEXsPalBCNgxCOqroSamLZf+kh7V1/5t
B/aaqxDsNrexhdxL+N9Qi9bI36EqCslxCOzr/47pZ+gEMdhsXMBrBva9uq0ftpebdQZhPMwjHliD
ESTLpJMaaQ7CsNiipTPtzL8F40xM+gjb99LusjXTIJVP/TVIEHxu1+nYTqN9JOPNPRP3WoFLzt8Y
hWAZREbc53rCjSPVUpat+028iWcyJ5v+AxdzbXOT7nT9v9ZVxoO/fs8+TRdX65clb26jyt9ZKxkV
VZHzNVRLW0MUzYh6r+U1Iyxqsl0yB1MDeTQOZBEMO4ZxIBoLynrV6OMasHExdQgpaYa7R6+dxXME
zrWclmJ8XmyaXETpVvk51IoefjKQJOQJ3DwMzUWQJtUEeaHqo+0jXjiV/rC9cM1AD0RdOK/v/Rr4
ThsiqULN/5UOm0EIc+D1Sg8ViDQmj8YY1Thhgsc/4T5nu5s2C6cGcIdqTAiewTQxHQavRB6S8i4E
Qb2DxYeFnH2IZXhb0H2nEKiNbmbGdDmwE0xcg4rZ42LSkMzUzYTb+KXV6P0dPsDSPqcdOfZgv5LP
z8WYs91+54Z0Fs9or1I11/fiUbGDkLwEUl9Eer/bUy4CMk389f4IFKZ7oalp9zp0z9qo9NxqxE01
fP4ZEaH9/YBw0UsXSCoEOWWL5VL4RP/1RP0GiuA3a+uBnh/we4kwOTT2tDHsYlOm9prXzE/In3jr
LxtCJfmxcdvLie9LifpByx3kR2RQh2A42rVkH7ykbXdjDArZ+G96xhcXCCs9LXCDpWmzkLlkNsWt
drTQrhIQriduHdCopwhtcd42AYcoFUt6NiiWg7V800QVV7GswdTaO9BaNwEtm0ZMHeH+eYzBHqtd
N5Fb4dyLGU79v3hI5R+2+iupXJdItKe8+NyNwYUXqrWS9J5Jv51YcvoQIJo/8ww5LJy3rDfkbS3R
15QCzEK0NJHkHcvulBoV/N4ftiBnmRO98xzifzykjhy1n7MsltxwJdMsABbiIWSt0u7ae/zA+ZbV
IElhaInKi8vUGmlceGMqpolfRw5WjS2VrI2UZCuO+Y8ydXsGedQJ7s4Vy2lIZPNDthPcGEFo9oKi
6AkSmxwZYjGmEDvRlmE12ZBO1rmy3oroIG6/NTlhCzJw3F8fOFy6yh+m/NApZb4pwrCxOcfynNel
a6ahjRRpi71PWSQSwWoOb/JEU2Iv/rExjJ4y3NzvF1+YEJy5akSruI6tDFnKnt3x1vutif61YQr+
KGCAQd8mgfDQlye7KYu2hnemDAQcEVGkmM4hN7GQmhXdNc0IKZbR/9c8cWIo+wHIuGPQa9r+rWvA
V4+U2yJKyFsZiNcghhYRQMAV6442gODhqnZWUgZ4O4FmuX7N51JiLgAjL07OhD0wWpQMEGIIjjqJ
hrwOdeYQK/JAd5Ii8gt/CreGTs/15ogpkrXmB4lwiFneIS1Npq1D3Q2jF7a88R+rfC4XA4LXBxCg
HEtgf1R3SOq1nWjeZ9/P0G0QwE1y1Lo6+Ukb1C/uVnph47ED3qJx7Q/K/SzzwREqDBs7Jlmq8AuF
WZwMCrXIpNV9iG1gcC2IsXtEI04dE1ogEi+jN44n/iyipZC+2+hrPtB1/4h4TY24YLsUvOrjaJrX
Fkj78YoCk+VKdBFUgcw69DRbX5nZsE7V3qirXAWMICTf9SZ3AVYH0lDweHjDqNty7XRQe29G8OAY
W3OvaeA3at3pFGzC4b8u8LEr6F9o1Ot7S/Lcp5FSwZ+3vVgk43yacrypOcNkdrIObbYUu4RisDgS
RpLBWWftL47B1ImxFP0U7OI9jbCNyPfcKNUVjAwiMlK9JQ6Hc1U5Z6A92Eb5aPNS2QtH+sEgouBm
VoZ3r/Wli3TgZEQAaTMK4x3AKihuCpUb4fyM3L1gHK2QpqNscGSgWyTDnAYnhGS6zTAYNOAPRGpC
R/hVrWKAlJ9jmsJjg29pm1obFIC+f8tYj44grQT9/INhtzlaYjIvuYoK8Ee5dGdGJ9xDLiVWT4pg
Vqyjld10R9GZrtLrxl3uYL01oT8YRy/H4PWPgt0cQxdhdvUgx7Btc+FAZf94DJtNRV2z3i2uXpIT
ABRHgb4Vn4ZXvUi3bJK9JmpGSfPaC6Eaf4pX8gQF5926GG8oM2ANNVVphyAzIB8+k2u+3i9FpoSa
htqfkpKXq4xSJMh6WDdzTBZF311QJbayoQRjn7MwHs/mGQq0oNhobtTurvnpep2LfKukmB5wVJW7
HFj8o+salZsvBr83vSRsztg6DFZF7Dmb9C5VKFT7pmAdYOoV5YzT/kGl6Xds7S6X/loNXfQTQevU
teLCVZkUulYYXZ9aNNcJmp9+GcYcBwHhUqRP7nBnauo5fVOPu78PAYbyCrD6/pkdMBD7Jsr6YtKX
AHz6Y9mj4I5FRKP27cB8WNa7WyJkH4cwLDpEU+D+cQaWF+/POLYbLwCBc1UkarXwvPZhNh+2PVne
VqR9s8exRT60rWoCwh50WEOvAUIfh9TEBuJBBgDM7g4Fm5fdITiwSFiXcLZzbP80IOtPUSQlcZgM
SuQ2iUyeV6kX5hqJqR4FUFamQ9ugkrhZKevTSOgPq9jfvP0egyA6hvUWYnYFyZf7HfFtI3rlstnM
OPJU5Va2+EsGBrr4U0Mvw4g8502aCjvvYPeQL0wkbg7T3E5HWUZvjitnqOaJlTd5HKY81gXB8obe
yv/K/S/ujaLqoeCwLNBGrDQFKYgyAF/TWhMuo+DApDiFSedN3YFzff30+G6SPLd4rTUq/VaU3m1F
Q867luho8YbMjO8SIOtV99Ovf/qZyHUrZo9vMg64VUjwY0EsymgqeZzXmv2rscvTHzKfQ1ySQY0e
bfBLL2SsZYVZ154MGI4SPoMIa8Ro3JXCYRKEPSlVua6eKcnXsfVYU1L4HTLa/K6ZGCLCmP8kRRRF
rG69VF+yP7lKzVN6X30p3eF1bbD3SEYVq2GHuiRUk5jU1rYORV2TSXH21p2m02D468aI7ljLVgRp
YEPw7b2cVgsiyYqjEKzJEOnAFrlC16xSgWAXEPo0RjiVsfIw5eVCjNOLyITXoEKjhnAyuqJkMkrM
32xwllW6zJlIckSjiY3RTCdQNgneGc4Dx0tMI636cfNzlAqDpqb3NW/2h7mbAFJ9uxR79205CpcK
TqTMd4gwPmKHZ3M0fDPCUXVYDb1vMSoe+dYH7/zkwsDoJXh4N/40K4G6jNHhn0adP0Vb1wqaFL5N
AhIwZFTp3r3VnXU3ELpT7QuOPlO69c3crnupfaXhIEGTAe1nNDkXb9/v0PjDsSA1BxHoRBo40t3p
Fp4/FWkNUidn3Pzk2RhwLx+4bV7QXxvEBtwvocg3pr4YDTZzC914fkTDEY+ut9HCYl4wbC3Kbf2k
aswxKnO0hA6godHgpfsszOtNqrOPHApW3rUcAgiQe8rJNB+iKngPBAaP458JYyVAzW6HaE/VQtay
vvAMF1NYa8kmm9CD56NojUP+/1enBHCgyIQ5lw5vpnjLe1g4VCTUNEdhTZpq6VWGVCnSFe5AKjR4
e+Pk1JQQiPwG7vRTncYiEY6s3Jk6PRsImbcSlssEuOV6fWRkiqyut63wGugkYHlRqH5xRS94vHcQ
BmMrYUzpEA32Lx+pL0fKclG5kRX6/Ri2RitwUqUa30eQu1uhgAGPlNVQjegAEZABCS2nlCipsctA
L40sJqEzW5b0tqADQb/azgTUdrgVx2sfBJd69TZbyRhqSnZaLJiItJ3Q2wg1tIfOsAjr71edTZtn
TxKbhcF3C7V/qeAQ2/agdmAuNxeTNWjrEGNlilYq0wzh47XdEhbODwqVT3HUHY5g6amdiIeaeiud
Cj+oOvViCLEbFs9UaGr3T/ujKN32TTHrs/TWUPKTkbVQ+ByKz/7wLqkdnASf6OvpToy+fcjr2u2m
NoLs3lY9uvk9CvsEHH7qY7JHmmVrOzyOKUB+XFz663u+eRXZkPM1NRrCNVGUfOTqnLOtJoOKi/td
LQYd1Xy8M7aOtbJSkLatC1mxta4U2Mf4YXdVOohrEP2AgqUIkZLgZ00EPoV5/euM+5unRMaL7OF3
NdKKkswAsrZaPjrJu4rZlUysHy2rbzfsQxiBXv9r6FN96F8TIUDcJc+gz158J6H0SzCzANPimIw8
Aacta5R77GqdactoD02FQFuhDJv+HaecKe4kynTp7nUKHb27qX8Am8CX8bMfdM5if1enk4gpvoiF
/vTupB9W6EkgVLeAH4jnM5YXzHJ61RhCD3Hw9JgioAVgFUirWu2qlw02PRucB6M4t8CpVH87NCyp
6Kq5ZSQ10dMIUUq12IEF3ZvTGD12vbo31lJqcaq0mj0MaAtGDq5Vl4QgICZlDK8WLl1Hoeu7Y8tk
grCEcaeq0Hi1ufyFH+bGiBm2MXM3NmT3sSx7kKfuwOAsU/LUzIYjYYrhaJ7jhciVplTf18C6GEQh
aQIo+jC9C5PMpRPQDXBtmEkrT/BAHMfvlSbCiHXBmWm0aHcTQFU4Eauhq6T24JpbDgycxpOYQKQe
2NGdwaqz2JE2984vKBnmY7PX0Oc4uSuCXdjHD6xiCmo0wnHoXXQ7YMNfGK9fCEJzHqc37aq2ve1p
jEGt5jSdEDFD2qwQIeSbKZfTh22m0NgPbWWSDWtbQMs+WEoJdrMX3RzIa42+qNS4BBNXl0FthSho
XAVnUi6QDAEDxuXrQBtpNbEta11BYr793Krdk6kC+tqHcMTDap1pPLsELpsAkbGLAikiL91zVz3g
Q1zwvOiL/6EVy6YqZE6RRSOPV35iUQFMEz+2V3L3bEADh+kj+ATExnpzaSTcMhd51QtFG6Jl3NYJ
Z3Jz0l94O+aGgsrdgaWSURQfntW9dDv8QjMCCEHSbq6rAixiqDDAkqmuUj4vkpmj638PDZWulctQ
JgVZasPLRb5359JZm9Q4i0Ad9oCmeGQbcBJIdF6jIEFykRBtWnKv/x5TbWJigfIl2NNqwfFXQr9l
n6ckI1z0zACaFD/yswp/9bwfRv4j3BdFtW6OU/d9m8o7itgAMVMVfdPx4juhtVwv4qccknBG1+3l
ux/KhgxmakaGcSTzCqvmAFIryIVMayoppd1N2car8Raerw2OTNbDc1/wYI4LWHyhroLv211mZoUz
zU1nTPGohPBj5s9vJSJM8OOJln/c8t8cAavXoecBfI9nr2hMoK/l5BWp3udUv63F5rTYnKQUOreK
pAuZwwhod8oEbEOIUjq4scGfb4o3fZwwkH9OtasOF7SGrWbErp+UJv6fDzacGPrWzIDStzKl93FP
UmlIZhSIYKTzD/1Fu+4Q2RPm4/JSRdFVRB+mx6GyhzemOLuxrh7QATkIgtPjYu73v5x2m9EgvPjo
el8GkjD51V59cmyyh79o+Zjc/e9NOMl2NVDNWE8CPxek9ZJPZAjm5uveLQq53m6TV2Rcq04MwmGn
EAzgTD6g7bt5xya8VOwmIiW7HjZ15oSFmmQ8RaoH45XzCb4194t+tyHEp3JBZpChqbNk1vmwwuTz
VLXwQrHYbYrN9z4EQV7GZPLtS36uQ34Pn+ywGBkm7V2uyQcCt37BIspVV1l2MZLyBcdwzHNvrvYj
nco56iE70KDZMqZRYMBd0zuPeLHkIENX69PCHAFAN1P5zSg873ozo3nxanefRY/HAX1xywFEiRg8
CTT1Cb2ln1qbHZPuOhSpHReEOgUcjSsHLCroBHsR9GKYchKRN2+JGlN9QHyg7yhAv/TfzBHUWoPO
q1iRSgV3kAx5ftIJ205C6oN58xMO2osQAB5dXVsSfuxftWBVs3NSA1oPqwBo9HgkUrPD5pRzYW5E
6oiHGLMVhmz64P7MRP/1PtjT2mEGi7vttpkVN6eJrnW4jyehAxjrXAKUX6P4WhWklsl0pMaj/6s1
Bm50taRu3fv/mA6jg3VMmelDh3qFMtnFRoxmjoLEvHGTvWs5DqR9W7wxw7iWmqlQdYAW3FmIhyAp
pj2E3g1YG1ysRnUpIBIImrYL88yZTzDCrDsg6oYP+re9ApbQeq2Ykgs2UBpp6+ZhJccLYw32iBCG
lVtzJ8iNQn1AAX1xHgm5GXtzpnV/+qVJg34+Q80jVX1SEHeV5NGxV9x2xkPlh3v6L9OWNKmwhp9v
TCpEWdS317sIyYlfWLFf0CEi3Oljzy2qEoUXZtFE1oDJq40K7c2JslYb8Z7dNSgMMxD5D5gB4yb4
8Y8xjWQ3AfVYFZS6aBYudGMjsa3Oi301K0afloi5HryAMndSfbk0JEDRcHAs8uSF30pcSML0A5Mz
0yCeIk9nZiC/v10CSzA3WweJysmXZjwl/cGSCJVP8gqtddWyNmDuk4ZDejoIFPw3sbfO6xd6tQV9
ESN9W/xH4JyOvSFzxyACNODugc2yHlvsEPx8QmtbfqzbhNgpYtUcj/BGzBBW5S4CYvPSsY6+hoEx
WmvLK6o59yPTzlM4F6s6z4uoEmQVXTgiD+PM3EODukZPr3dJkjlykPbTCAfGNIVaXp2wk6vte/XB
ZTnCtbJcX+nQcUOYIiIbhFP70KW2Aomm/1q/c10gSEuSbVlMIPMVFdFehox0wJb6mJCjjMAPWl7I
xYIJlIokydfW/kHrmiSslzLfeaz7mnnMXm3LIarWt882121iu9L8Lj6CbHkd27y45C8eRcdwRbDn
D/Qz2pC2/miLDxR9xCjOE7lZYo66iNH54SJ7cX0ETuLuRpztvXn9G/gcqRijjrXKBpyIzKSCjXGS
o6bOhg/f+Mzh8TEwM8ZelqS9JWvc1DeziKpIPmWavVpQbdT8YRV686qBHDDm9nvYyg8Ddfa3v9/I
3kdAyvu0TXKsfdyJ3ObCZSxTHjxvH9ey4GBdOK5RM2zdsn8D6MBjxbZMZdKStgh4uKwj3na+vtEJ
ev1ARpGrNayCv705XE7aS0K9uqIkFCxVSRUlKvkEjECr2atT8ulkoKJ7zQklM28PNSM6c2j2ZD4a
GrNY6ZYM5Uzp3Ffg/rL33vcbbeB98GZxs3td8kAi8F5tkNvGvRyXc/jk2kKg7OiFDyJILsZBOFLN
xjKHFNU5YHVN9RHUSAMCdgIJHXw0LLFx7k6kzfLLny6J1wXN3p975qNkHTmFld/GfaWk+2acIdWm
n1718IUJgkKwacwHbqB7pQUT45FwwiBB3XcWVn9YJl+KZ8+x30h37ZJyY4X8QOEtTZYYnpTO2zOM
2XESPbFlRhbI/jLcBBYYI1vpnF3GW7OXFwSa8KAfoaTkQTa58SxO1JH4nzGPfKuXr6OjmgUes+J1
/lH6AEHe3nBYz2UEcInyCdedI3Yjj+jf5WaZIX8xaQ+cUu0wKZiBIIDdnHAKxdZF4l9R+/oFiy/4
obQlTEyGTGK+nV7FAKytvnoLLGaUhY3UfaVWSi/jKPwQ15gsO5LpcPxY68xEg0p1sltRslIoOwUx
zZdw+LnBMNffRJFnYeARwOwrsearRSz8+JRuY6wlEnMr1kcA7suICzkV6T9Fnfn0qRK6K87vuK4A
A1uEpRYOrMEvpsqk4GJaIvtGW15xqDLfQkqsLTXjX8aF/TCGAKg7wgFjwrV+J6ZHrLsm85x5sBTv
SryZpXL01aoyYmZyRvd8MzATVtxotyUycUoDSYNiZ1ovBI/qzrePflBqK6JXy+JtHyEzoqctO7JZ
11DBpPGZRq8XWPHLUQh+C7owRLt5/l0PKWgdBQC3LskM2UJVG3oiykNa7b5bf9l9ol3PYyYfk1ZD
oss7lV/neCZLEaBuOAMnwRs3B5LtXymoqXw4zn6lryGU0qSHQm57UPkjA1rUg+9ftDosoVM94poW
4jJlmFkS4w10ru1gv4G3v9NkJ0UM8RyCvrJsml5T06Op7J4IWLn05oJaLtqjxeWWdvNtRApDuGEb
1AIVMXrWOkvy1Vg8TbKsT2XVa+3LAwc3bFGWg3WEu4MILp80FT6TkLkjS0hUFv5guS8UShlH1Fyf
Ci9dSnj0XXot9LmwIjEQXoDH/h3yoKOxoraIdqyFOtT703BNn2L4556yx5vtwPIh0NclvDSJcR3P
v7cXznGLpvOhXLDfiOzxinVEmgT2xDrFsxM1smYJiU6CCuWehUWRfWRqxQGQb9qR2/yWw88sIO0P
Qj87nWlNVKYpI8O+gO5G1BEPalUKaH2tVs/1+uMXGnQR9ABTd2HCL2w2L2U0pPHDL4uQEu5MR1Hc
fdiDfmkSn5vfcAUf0dtUFXPB3mKYjMMtfJok3QkFtt/E47hk8e9MqeY61inZGcHeQrtxA5fPyK7B
mnUg5XcBSScpeAFwhwBLWQnKh3X9Cqg18s8mvjenzDVZK7fQp0kQC2qW2prXTptwuHEY9dVZOkTw
bh979Wsgd+MN9PvYFwspyYW1SPfI0Df+m+deKFOArmqUQ4bFhe1AMHBXKtOIktUYbQPlTavqvnSO
8k/OxMMlxeZPMa+tgksier16cl1MUyqYI/Aiu+SB5WPqVOOBs2/Myf3jAYW5AlezKxR7XGM46sNZ
KAk2Wk09lp2ZKj0FZK5HT6z2nmeyVSyHOtpd+R0qnjaLqgvA7Bm4m2lMMozlS2OEVU7hcvWSdzGX
uFBuq4mqk+mgeM5shXXhWk2haenR7B92hxYsKq7x+DkmgBxhGYA3DwdHrzs+6sCb91SXAvFd66TH
we45UoxJ6ZjfWPeTTFsOWYaik+1htYNRCH923wLfdeiZd4A7oEoMFDmKi1nrMntg31iFog/EE7ow
0BYrf1fxa/SQWMUwPQ36PdE5A+fU58qEE94eUUxM5SMrdfJgwHLD9SiMTCegN3oXP2nSCGqwqgYq
F8jfNjux2XXjALJ27pXLZ7/sHkzeYYBqUwpcy7VIkj+w42ruzOHmrCr7WYOw4Q1nEidV8/n1aN8u
LOc7XwfWCRgjjEgSTfA40QX56Xtd/OdQcBNXJllRPJEzeN9DNMClPWPpBShBSe7XyrgYWFz1x8jD
bfiuuzY1HIt9U27APG+Wn230tdi7bto5EBcE42Jsgd4LUKUdX2trNYWP1JQ6M8mXjrAPPb5hgmAE
xZi8bvsw0A+kO3cQSQLTsA64tOerJFttZFI4gc7Ca2v1lZtyX18iRzwIuhVCmmD6z3+xaTkcHnKL
qNCZd95mV9BRdZDcm/euL0MVwM5BACYcuTx/WuXXcfSzv7R+EwQPfSO8gjKPa6uthFhXGGkUbOLW
9gpfO1C6PNstzhCEcYCIiFd33ZF1p/ZhsqeMXuNRavfJxGqI6vMRrsMo+wX0omKxZeJUogDbkcVO
ZXnRYXmC6ndbS4ktu4JJU/N/sMOfLrCEiFo6W6OyXTvLyfpSfJg5qKOmWMKPjsGeYVDlDw1kVacg
VMhaJBQcOBDlPvrjQJfRMXRzV173+J6RkQcWJPcvt1mKq/rL598skqDY43hfyxXZhodqWYgEoJQw
y6OnZAE80GZMz0nKdVRee6+ZeZt3j3Tzr1zAdm+gXoEDbj8xoY/OSavOI1gP79HxAuK8HfNbNmlX
DfmHP9G7cRhQ/+XRmqEcwNpZm9F4NQk8+Hvv/04Rv/rHp1UUHq78VPjpUgvx2EAXiRaqfRrqqm7M
iJ4vxe/kqxOM8hvV0plg9jIpGfekYi/ImUab0TV2ZnxtbGIenL8tN/Y5/vtN1SYSpaI0+qp2ssiU
c13ucGh4GEJXas+Cc/FB/6MGW8zVrzoBabxf3OHm8EGiVVrb/ks/1mEn3uIxd5baDsLUqXEdV99g
USVGv78M4UOLjfX/nkI/Wys+KzyehidLl0o59VGtuh4LXlgXeWqRtMRCA3JH/OHefeXz4ER/QDbl
CDinAF224a1Ux27W1zlqZjekTxoD9p+YxAbmyVT0m1mwurFkTSKtOQOav1XmyyUVJUmEoLZ9V7P8
gUcru4RMHftRSXoV3ooUaFmpvjJlvyZe2hUS23Cv9KvtQj64kkr9qhGJ3UukruwaDR7FineyGMOM
ird6lKUydW/lwGHXwmj7m1RUcIat1hkGsRnaGIR79pbJmDqE5aKSRYpn8l7vu+RYGN2ab317qubV
BaCD+prqTGrSf+8oKCMh9MOt2OIDvWMoRfipaPzhYcu8fLAN6WapO+EKasg9ZxnAA4bDYIZieB/Y
HL9mh/nlsnpQNs7g/5q3lY2ik7ZLci7sInfM6wb4XgnxgzlL6Dz8hUP7QTGR7RuUvEjiP8jxq/Pi
MnL6aHhNpIdmaitLGUkjcgJuJW2BwULzthapMAri8rYFAGFdX9nKVetYcTSPAwdcw0p9hFw6X5za
Lkj2yhYBU8kqwK537mjg8C+2eQx9uFxWPPg7/m82p5lKhIkdeSoB8x3KA5n1P/3c0gaDd4gpHJ+2
fzHdxh9SuDAp1OUVORBS83db9RCDHzK8LtyVXWAfF/fNRMo+38rPi1xNnPZtqDLw7yXdHIcz2tds
/KxdYC75eNTxvU1gPzmWa1v1+M2qrto+JCNzkRTIMZd2kjzgyZWfvv3vmnD58R9pFGRuH3EKTSbW
W2lmhOyAKN9S+4riPMrt1fdeeAHK4SVzbqYQNIkEdmuLohx4a1w5QGrqMFc6IRXBf5OJMFOglWrd
oJbsvanNYVJL3oYxFLRRPpoZZPoZ+ppw7sz6GhuPlO97ifO3Mlv/a15Ktp6gzOgdoVPjEQkw0k4f
GLfM2mAyaLJkiQZd8lYIUlrbXpMrO7OqxVBpdejoBHGHk+qA8OgzEbEafM1PqHwhzdLxOjllKfR7
lZoXK459Qw38dUOxhNsCE97Pc64epCKhu8vDwbKGWSfAB7G4SV46uez3Yv8JVsyT8p3AOahG2TrS
udoPw4WXJPdcLkkzua2CJAGt6l7hFeErTMRyqbyA7jAW4RIN0kGV5Ab6G0bxOzghYeC2/gaEbpxm
GuuhUquFB5R0JCza6anoGtsE+G4Bq293o/mMXZpYqZNnIEKQTd9HifM+Nn4h88a/jNZKjO1sh+KX
Jl9nKW3mlVWuklcLng4XZXMJgiJcNxo59o257TQujgF5HNQNFrEEj/tT2G2pkf/C9areiNhxdSuN
ZZe8VBEc3422Mw/xem6PUpuMS2CDaea1Jn6hiWRK/j6XrxBcFV5UyNoZNO5XSVYHfwAI++0HT8ch
sXtuxqqKWlVCI6HiHcauo9A9EcRaVfB/evT98W5duTNLalwaVfnMxPN5IlzrOmiM34NAE6tk5wVr
JVlag6Og7QFPe8PjRs9D5uZGP3r/W0tnC9X6KMmGxpOJmsk1TlsWWNrlVgicvUlT4LHiRXigwJpe
jeN56h9dAlVciuLcwy7I/yLrp07KeJ7R5TY1zpYxUdI1C9loQDvu/jVoA6Fv9PcbMPENcKbUFu7y
/gU7/aRXDqXW3cFPG3OpBQwTBE98snXT/P2IWDXfcB2TTyrY3MVHxRwyoWWIdD/QwzoEftHHFlNn
LCjGaE497E6yLkKumFjpVZdDtocBpDxTVuXbJZHBhwMikn1BYbLp8Y5kIQgntMJ+6bOM6pYb3/1J
kWFN9jyJ69C5swA9Q3Hwonb5czj1t6SHWvflyTUHCnG2UOt26ZDFr622t8kKAF8YBwBuIcxErX8j
8CyDqJwOTdWRJB3kNpwsss4mCpUe2798a1A5CrMr2QLpnoAbmMBH4uWia5eo1D0eb/HM3RrHqXNh
5HdXEiNVHfAvR+eWjZmhtTEsc9Op7T0fSzQ/xN4aauJLMpzrbdoHWb5fnMUNm/qKjFXJJMBxTFDn
7G6ExXNTZctwJ3jMw4jQlZSIRN5XmqQNvQgh2uTeFx7IqytiD8iM3wGJPes1j3RfC9mKfSjNcoiF
mlFdjx92foD8Q9l3t+eEBEaxcLVxiSB51kkxhOMYU3EQPx/K6dg4KsRRlWBIxkRKYwq9JzYm2v8N
x3S85+7MfsOoiF7k+9rtBY86TghHZbm9jbeLh4a/9tV9D/vaTpKA/koL8pVRA9wmQh0U3p1Z78Ba
sdAQj2jmh2ebjjV7VSPcpSUFpqv1S7MAzudqGBgzpRq/XKxc8F4dRj4weWiYQ9m822oB0TbSi8Ti
zhXu8nR9/xZ1UMBarQM44fcB1aSUvkG6OXxIV6f9eMnrezj52jq/YESgyjhbCGHYvbRv4CateuqI
nQ6vcKweQCocEc/1DDfNdRK9lWaK2SMI0nedUX6k4hhmfz43FUV9bTYhf7awTWIoo06ea/mtPgX6
BdzmWZ8dTaAKTjWq+9UcaAqLme2/Ty53xBdYK7zJT7LievK2Ko8hT444MaxrYgP3yq1miH3rHV04
ux7DMVYCDhHEgPSChvFbHts6GYukXHzagAE2sJsYQ79oDyCAHpMdmvS1FlfQMrP6Lu4ggEIPYeuK
oKZAJ5IGNGdwtNNvOAWrbCgHmYPUALlIJeh1qX0JRsRowPCj1WTTU7tcWIb5QirjpJULalDI5nwf
LhPCK4Wrv6fdP7jjCa14Z3yA3yQQbvl0R9NtkXQQcqQRPrrNGS+BAiqjitk04p3aL5IJuzh6HTTq
gBDfLFumfm4ymdE49nVx29A3egfmz1RgXbIkEKKELVIDhuNY/LDo8QU+rT0jQKKAMacqn4DF6zFQ
UpohB5kZfPdC3y8EkEyWsehS7UyE34YTbpjmGggiUrLctENsfmmpcXIDKqmjBrgk2LZ8pi7wSG8C
RDwRHjlauU3s+jy+LTqpmVzx1mWlMN3mgHK+++0lYvICUf0CvCFipJOAWI07F0XXWYGOb9cTs1CG
i6aEjJ7adSVSkNR+Qm7LVTTDNymJZjJMvi8Ghig2qr+diuopQqm9JigggWaQo5/lVxfkbgMfp+gE
Q/1mItc16PxnqijZuftdMKI2hRXlxEe4CqFOzp+GsZTvH3xIOJ0Sv3I92QOssvxbq61mQD5oPgha
V8seoUYKD2IDKuYObvX/6a8e/aUYNJ7Go4Vyw8SBTmN1QXjfrDGG2jD4OenoJtp11Y6X+7D86POx
abqToyxAnXx6FwvjIw0bSO+gN1NtoIXEejjheFefbs5sKV0SNR3G9ubx1CG+yxci3Ak1rr8VI/PJ
J1DE+B+gDlUojdEDg7KKETObwS90KimxskEQ0NwF715JBecPg3jRZK7yfDtY31GxKYrpyE8db6Vx
mWH2qYhqEmEEo+qJ1yca2Myu5W2eOoFaxdGCwy3nLRAfqJhsaVUsxPnK4Ls3DwZdDP94XtlqozGd
rE9HbWEsNmSaplwcfOvhsScrOz81+YFemG4u5j4055KOgIVHmCBq42d/rpmj9JBkcgPrq+yV+djp
PJSho37c4Sz/tvAZb1rVWfwV+1FG51/bcMQR+liko8g+lH97xsbMAtqaVcvKMgKGxWpUWWt8UPOl
LG6TjiBfN55AuacRPcrqGvhSltWH83aqcMGPNjcgwaQjo5r1yQjjpy99F9MKo2IOzVBZyC1W2d7F
D+hdONH12eojPzYJtno21VzzDFlei3r1y+khyHYJuhNLXQibCd4OawepcO1dj5tfr7XIpHpzsCtE
e4Y9Yp0TQK6CmcMU0MKgz7yaKlCzgO8N4C1vHP8uPuJzc0uYxcnMvc7OxonD7KSDkRqYtNvJ755p
Kp5O1+simwWK8FHfJ16ZRqzd4hpYIARZlGFuF7jYLvA7B4JRmF7+2v7ewhXC1EsMlGn73F3V9wTF
5kze6yU7SZwuTRTGtuvIJqD2vY+bl6TfTkO0rxsYk0AzILbq/qBOU1Zb49428PXRxwkbZFhyPjEu
shLkbl2o2Acio9IwiPyzgjlKFnWs+VDgBbARDdewl/WyYUXwZ2n6g0twcxLiNCxyJd7FdDzE6OdZ
W36W9wS9Jn1159g51MGpBmriHunh5gLPQYKPgIEqcQcyAHjXrWNWUEbVld9KIvSHpdI8KMzB09kv
EWwIIjKqhP8yZHbroVcSqMch/iOG3EijWrOAByLVFd8ZqsnrSKWQGKB8X1UWPtNfRBZoszwgnfai
hfH0N0V824NVXwbfQ1sKUjKn1lTZwi2tWUVrrVZnyoaS6r+INsy2jBdVEe683TC4CihYRE4es1V7
0x3mteQBstEV/wnZBPKOQOxgQ64X09Ot3zlcynyP0ZbfIT5DWMFfHhtpbOPpjbJBNQFWn6TLTL3e
0pC2ptheDQswcw9IwAVDtHC5b8AxpzmXhv5GOM5dfLLLAwEB/2AyyvIF7hPnXkiSx1HnM4oM+2tg
r3eBZ6VD5eDO8BVt+oBqKlC0HIMNyoTDMVaX5PmEzerCuPgnC/1axUFqWRhgtIbu/w5qlBJc9ibE
7T8tmzFs2yRm52ztaMsymFtol7duQTFbKeDD/8We/H2VMVYapz8DizE88709jprKzDNwMSbBCfnn
iU4JZojm+efC/qhbHfAYWhxOHT9mTpt2cUgDLQsS9JouUh6+rIaWhp+szuPyxXJUH3Y0xQ+myYOa
i6+vwTSD7g9ftoszEHQPUeG7FCidwXb2ZyZnkHhTME/ODb7yRbvtUUBZd3aNXyxuh8gvpPmcY0iT
EeU7tENAUd1mO8bJCAZPjxcV3+5vODe9ZInfX44/J6cDxcjXAvcGvdpJ0lR2YbhB7P/5oPrHp905
/XpHzPF00yDQmtVBg7FIcP8gq4j4NHF9eKhBdIlNK0AEH3kLWl6gMYEQDahk+kt79fpTzcNYUjOh
73Hl8pkSkzAvD6Qx+unbr9jGPsU98NeqzUNKputuIbS9FlXdNxoAdI+kgj1YB9pILeepVx0SxYVx
BoW8ETTdEQi4nyiq0OFblefOolKMGg12Is8iGFUhyX2XbqqNt3sfXhtSFsB0nszTAxWguzUvfrOY
KaLr7UM1U6Fa55yjVFZC1KpxJ8zr9xdzgTXmFWyll9pTxWxXbhfbntYJ950DE6oMQIiYIqjFVECy
HxM+/ziFIyoP7gfzegYnudZCgocsK6lNCzgIOGjK7Vu0gCCtVCAM8ReApwxqXIWIyoIY279ZoXuq
/Iz5rNdnWq/F+DhCPlUHH13wYSvPuN6R1Rk9wxLmlHRzPjGbFzlpugva4bknOXh8260WyK2kOPOw
s6zdFWR37P1KXj7PVrQHGwlR0yj/rOrva8y6jcJpj+5s6yxHQBkWF6S6iplIz30TfOMMoD6M9Uw5
L0cAEnpdfeNSdgz87Y++ybj4ElY7JFWDFxCaB4oQzKI5tN/WiO+P/lAOmd0r5jzXmKEFTd4askaI
C1NJYG9Mr9trcnMecoJgQzZJ9qmMO+mkzQ/kf3G/pAbaLA8esqraARvGgDA8KOPLVe63+K3N27SO
OMF5vF+EJ2qtVF0lc7d9tAsyCQ0vy2M1W0L2I9qKznspSlRTzNWsXkFoiIQs1iqxFOdlK4zCatFf
iOkgytpDDIsGEyVF8TzB0lHNAuUA5PtweuIkyiWTpE2WbLFcDHIy79DnmzuncFF4gMcfU2CslJ1p
/4+XitbcCkfGGx2DFeRFf8q2k5JEby0C2VNLhJE2deqv0z7bUIeQYWjLyy5Ca+CakV+DlROw+UsR
wOKz4CTg3FBVuaxWWdkE3za3c9wI0bmal15DuY/kfyYa59AaFdp15u31Zuzfo8rflkCgDH2m7ktQ
STsxvZm2hNYYMqMVkueUS8Ce9QCCwLKMwPqdjTmL37B0g3ocG+H2Q89HLaBmA3qXEuhpu/SnZy5e
eEQj756N4pvQ/X6OB1CSCebEVz8PQDlNKNjGKj3HZOZO26MUPanKrIEkLhGxoqaJwMPJFdceVDl4
lylmaxVri1Xzq8w2f6Ya4mLs0mcZmrVcyQB8Y5zVTQO2PiOVMkCFAC/nBauqbN6+CBsjNXaYbmDc
hVeRf8/yofTvS3T5kwACRDC8nwkJjlYk5VsyBJhVQtiGK02Dj3R/Q6cSXKaNPI0CLfvJ8rOz+Lsn
CPUPJpicHcJ/qrUZFG23KLD0Et0I8uvZutdXw995+/YkFKZ1+ZhURQjynKpR7up7ZYaoILdIju5+
tv6qAanFXUCcUy4x4DRnMsbEJTwm7qauDgLnlTxcYaF8iWhEKfqWL5Ccivq+srYluxaUMXLSj8M8
jJHhhz1vCmjhebyWcxWu/VzFPTMY80mQsRISCWaYYth6hHSyv53EBRYgewBftQXQfMFgG3JTe6mN
dpSGYvitDRn/NN4hYWppIsFQMbi07lnJ/z5hiiRwRanxhQoBF9rXTHAmFK2OS/Jn+s4hifrxRr8C
47cTqsFZtGwFevqwz0CN4yxEYrwUH/Df5ENTrBkd+f22iiYf600rcuCqosvhg2Be6pcAI9mZNK//
TzYS9Yox9V830/HbJJ7mfXQuGSuM1qwdeSn4gV1qIvFcBZXwuHAWPc8N+KZpXFutefgzFRFuY+Qr
oyJCemsLXbK0fNwDJn5Ha5cSTySTNH02NQwKBtMDW3Z+ybBizbQM4PUXjBtxWq6dgajISrTO8o28
Bz5wN4kIUazZ/2qPU7G4sgHvFg2o9lKnzC4exI9reKdamkJOvI2rNb0TZSB+zKNgzb6K3haoTkpk
Hzn6sh8pfXBX6oBK5PT9PlzPHX0zFVgJj34n32YyuLsT1XKK3CKBU8W54nCuJtBOcbbg52Bz0Upa
B4z95T/+ZubVWRO0j0ntRWsmp1t98ksjOkVsbIFpHRHUmrYEMrTdoG4yFSucGutfqndeh55Zq81q
IfYvKPLf08BHlB2Wb+iFdsSzBxmvD0CxbDzMrwvnHr8TKqhvDkxHeO99Ap9xxP/fcNKv5OESoR9u
E9QXvICznJW5viiubizp0KYalg3gd/set6+8Gre60JEL7J2cG9K/X1rP8l6O1BtSrl6JYDfSynsF
ONtp9Yz3e0OmJrP39CqzzR83I56g0UK1WnTRg1AW0BtogPdGbUz7IKFOGt2IQUW+U0H6R+QlYrnJ
4vdh3AdPPLkeILXjhH3tvOyzoMti1NkvndnrINiMGSWMeIHGlupNlHq6tEcTeSGXl7ryD1+VHz9Z
3oVRUk7FOq7UM6I9bCD73sFDqPUQ4bxu4yDe6L42rwjtULSy7Gj8gPeAzTySJl108fdtE9sTXwPa
e10J++zzc3OOYxc3SS8CXxyiPyx1EKkPU/JQHa2Orcg34xNyhNElB59bjjtDOGByXK+nfW9JdWii
JMCb7zcqKOwyoVwoCGAUEmPHVCRa6wHvMc8qQlLiY+x+kXoeTeJllO+z2eUzk9Fdkz/UBM+Tld1b
lV/1oXHNZC1JO/hgLLh/PLu0LA+BDX5NiPX0TVpWquBrGpmyroRbNJWepj1AOSJRhpVYBUwYGHPN
mKoHr8base7HhFmlcyH+0ODnf0K3RYO0HmQA89ybXbNLeYfY5/MGCQ04pKAJd0CuWD8Gzxn6pQJn
hUufax8J0dqeyGq278gHHzRVLOhRMMsD3kZyANw/oixDKJhkNwEA90yOR+kZh3p0fM59y96c0lTA
h8Tn3c2/iaj0QsKYASpyz6XDLQcJCmBw3VlEhcCkSXwKN5EvO3+4wiI7Ea8TgADC+NGuuc46kRUP
hPnDg63n1FFMptzt1FyNN9mSevq3eTTC4/qQ75QrJ7W4d/ut5M+OV2fYyFgNmqSbxH8Leiph0EDo
uL2DOC074XpgL2IwoKLR7xrtydgZJTOQxTzY9R5+h8STOnMA8VJolL5PUTGdGQrXBQVz0UeV7yKX
975ZFt1HIBr1r/WiggVxqLXDE7v1lwyVaRcQd3P+SVPXVDy7AWDF2BEz7g4cH5CZxHqqERgtZ3Cs
cSH8/iFUHozD7qFrTGN71poqAaR8OVFSBT943OEeXNsT7PcuqJROKEptT421tt7aIJ4KtjlpQwjO
D31fnJQUXKFWMLi8X2B/RCoquTUiMIeucWrZfW5vp/yEUmfSfjM4vi9GLNp21eZoeGR+EQNMbOI/
4q0rnM/fvCWCkP5d4V8GK4BVbv3dNgxz+j4zCwGOfGlCAjKTopXPNwSKGzzSH7/oEW3NN6xJn3rM
xwLVtPzwORSAP2YcrDB+TThSwIw7TFokB8l8+AaACFAMJ/5KxRV9+Om9Z5hZ2mngg2uT9K/8Tp3B
Z9Kpoh9aSjM0IHLTc2mhCkv8b24SYXPzEL+lXlqXWE3K1ivF6zKuzNYzgqKwBMlNFpKESYYeWnHE
Js22+6ndJ5fMr0MpMsM9FjHnPC+UGM76HuhaoNHNPlCAVZRGfFYBSEf6LzYhVWdZM1AoerBjOmro
LVpCQZFGe4V+kQp0hK6D/q6xTDnvpnUPkNMHGqLRwPNbDFYRPSO23m32WdA727JJ2ftRihR/ypKz
WL23O0PH4cT+MRVoeU+A5kjZRczmAC/l/DbvbBgbDpCQe+hQxno7j7qZ3TPnj1yvseM2Z+MMzhYI
TVcm31CfkIXaSIDuuYcDLoDDZTQ2/j9sXPwKEpjJkW4CikdaDucKKJ2rORxhM7FeUcocCG2bfAFc
8PvMrQ/B0B1e15YuPloxFJ6tCKgpUECEKOEtCTKP4koo2IPRVQyxx+jYTWYTSMzKGvBX3qL5AK3v
s0vbM2QsHzjZU44bGL+Rm3M6m3kLbOjKpzgqrmfgZI6kgmD4cwKh/p56saxtHe4vAdC81noYPOsS
P2Bjd48DYJ/hZe+6NxTU99011NX8fnJgm8F2grl65VUaRSKj3JYC1nK7EDMdGFA0846bN904AsS5
5kSS6yR5g67AkxwlbnFDvXT0tqw3uIwopeirhkmPmjw9kjyOsCGYU9LFwhvb+7LeU0M0xOWGRBkv
6O4B9C6P5Lt0dG3RHK+Ohq4ePSJ6Kc6x3INVGaP/DBjZBn2Nmc2kYgiXkEjXfSd8w2kmYYjAGQ+T
3GnUahCX29CRxzU3IalYd800llHG/sUuLB2D/Orrsa+b9CK4LFhYOyP2DUiIyujTWaLANwjC7R9Y
m3UsHwSKX6ZZts5DDNOgIytSB9eCDKRTdNwEbCAjvf7rtoDrZbpbUFF+AylAj8+AoMOCbzUJR6TY
wdgd+TmFylIIscW+ay0EjQkYzOWCrCQYBs4BewblK45wuX01SgLUTqDyPUwYk2KOThW0FzHv7YZr
0eRk93KV1lMchCf4lAiJsu9PiVQ3MN/jAaig+X542faYOMvYtw4n5LKvInWzNdXgC7kKyihAlXZI
DEaQXL2HSh2lArcv0dMHSTn07QKuET8PubVnaNVgrlPGSAGuc6l29FzxsYWAynj/bs5twlQ4iNIf
mnfLZu1jLGC8iwOd5aJ8BgToeWExGbtEXJdTvzTDmq1P6xis2yocnBnaLwIpHEQaUIR0BVqA4a2I
pllH3/PXyMt4Yqp3O2UTkT0PvcqfcmDmRj6BCykl2TP1PXVwjAqAa7BYgH3loWnKWAz36Sg3CRaW
BEmFuqNtSfhWkmQED0SwK0vXT0z/EbpLtyPr/5kGj0Dj06K3Lty+4ThHfeydE2Zx0E+4P3DIS5Z4
Rhqi8o9rsVcsgXndToLi3Q2a4fDBjATDG10kImON4ecCoGMCy7HswDSVHkHVwCjj2Q7X0m7ZGX/n
3ykqvYvdl7KZIRoTHUVcNlOZMH10seCiXW7DkOO37OrdEXHbm9tabcUzqVJql71xRBRVXNbwbku7
q4FSV3liGAclsP9BLMY99sR3B6fnaRukRXkv3HgqI0GmIy2H+tcWB5PfzQ06ijPHvr+AKmMIJj24
u4ftsiqUM7i9m+hqG2ZJ2gtDeZaHcPjS5pg0//Qm3bf/sI3fbJSIl63gwMKR7eigt4KPvw+BXpRV
zoR9kKUqz4kHZC2KyPytKgwbZrluNoIxbn50wH5PhnxX2UtNdim74GItm5XufDTNYozyQ8Xg6zKg
pi1y1/5LpiZPwHv8wOz0OwlHuBOsCUVKY2FSM0fqVpCgEgTl+6qAfB9fCyTLS4GyFfmnKdCpQSFV
38tMOs5ysTvBCze+m2lYZiwy7PQQ5GfCgF/5BSbkkde2Vu5ZYxxdeyjpkGF088UYz1o4Tsa20tTX
UhA5asA1fyrz+BsUY+U4GzDHOODjQM/Mc++Pm2S0e4rZSHGlbIwJxHQJ3Q6tpsGjkXkP3OLDk2C+
1fG0WNqWnKJdUKYHg9Kx66ZQ7Vs2An+fpwKjNTH2+9oOTlammCLiTVMUCPvoke5ulg1oxewg3eSE
UUU7/xlnVFOjyMnwr1wCOl2lfgFAxiOZNO/Vo+LWKeweU6MkLiIb4GoXrG+BaqK6Z41LfxH54T56
2A5CkleTsnhiKo8f8hss+ZmQw5RZ3/pUzLnE9SFg+AQ9qfjab+TcZWCB/LS8lM3fah5vZ0nLH9ff
O1G2fJjoC6fYomD2ycitUyUYDikMsiZ5Rtb6Ncvdyjs/nOIx+17T8wP6cSSw83Sv53WUR9BmX9N6
cKrV0t0aienj950yW5Y194xh7dnEoA+NsbsLXkVu/RtemiU9JvKpoYv5aKOVXZDetkql6T1U9ab9
3hVcGm0TxNQ9ddAo5WuJyFDJm+MptA1I42VjvUYbxYtbAec8AFBBsNCaUy5ticEhWTfLLG3sBbXa
C5+HHDPsYhn1Fx/P22ydB2/Rk317n6NBmcT2dxWf7PdWypF3XSlScQDKI/t4FTIkYJUEQ04lI5Rk
c52dJmEC3Vy0j06UMyU7EnjyOBxzvv7Pr/Tlxc0uOqBUhL5FIRRZYoFM0oWSOEB/jGzZoSncM9MU
sJWYrjuXk+YGHaTE77s1r2dl20GgOrfk2khncZ6GpBYaO0Vg/YpVm3WS/x5LK4YqfNn69AKo90b/
WFJXzsKOAm/a981VLCfMvGsbqdfC6Muiao2d76+AnyWoMt2XZJhgP3S2T7+1X7Pet2aj2fB+BuWM
a61LUg/7TeWmhW3q3HHltEuQAuLUhC9povYYwPmEIdn2r/PBDN5Zl5tRW4XqIwQkw4VUc0YqRMpA
NyleDUinVCKX+MeGCAB7oiSVIoBrHJffH+2Ht1WUcgKvyY7r8Nh6gRZRt1b8pcjWxnEoSLSSpK6C
laijXsfrigYUGH+qBqbvUqeYCZNbDKDQQZa2TZDo0lFU9Nh1L/3M3Wwym7EwFmqaLwqjcxYcqBhz
5xMq7o4e7qYjLt3qNuYbpNuxLtYmqoAB90mjg2J/Q5uyGDhxTOwOJHt5B176HgOJlyp3h+jUVCc1
P0iS4Aw0gM3G9KO8VSycClLVhakRW9Qg95FUCWcjVBuVC4Cu8HUu9JzwINty6euOn8ku9wEOvIIJ
ilo7N0PEzHWSk1O5obPr414pDyLLojQb/QKEoctrwNEyGcDb8ULsolqJm/Zf7YtX7YUPZvlAxJHP
RpaOPGRPmqQVfX46UBveZSPzkBd3UXpS4jhDYDEaYG1sjQO7rrUCPfLBzx2yVCFn01Wc0pzVVMrY
nYeGsLrCaywxOfEdq12ShPRpB4sAGeWDnX0ikmYEuAi3DikQFhd6+3HYBcddKb1K05qTqYSg4JW8
LcpPfpjuHGTI0FXE3utaMJS6hSi6oPSgWndxlbjEE88280zzG5qE7nAt7biUarELQSwW57a9j8CL
FdejfgiI6MSH+RIKBCEm+SbXkNQGMaZE4KttboVO5cIZ0BYn9GtCcfsK+LUNX0TSMOosK++oyJsc
WuMa5TD1zfNdXlJFk1ZJaAHRNPE3Nv6jakmY4cOM57KipU9EhcUoy/JOa2HOZMnZnkJyQoBQ4UsN
5/0u8sy0/NupoQLEn5l2KH09D+OddlTciWTDORB3+ZyeRc5f5n/t2S8Ps7VkzNPbjggWCKW/Mf0C
OatmbkmmYH9aaqMsIdV4Al6KD8ge6yUR3PIQGoQKZocipvQT9TYNoUQf5uXwy+A9Ue7a1xkQUMOS
busVPxxG7CTk9UtQSOisK5awWhqwgU+7bCBJ2iuL3exUFpOE3CTv3+CMSLsepb/UnqO54BJZNzi/
EDMYO3oWi7Ull+CSr59MwzkHCAcTcImVYnW7b/p5X3g0KKwRsbPDtWiG8ntZPFTS1Q71lqozQtuA
YFf11l4xO2ICe102ykHgddyZNTqVPzh2FRz/rS3Q5ZiioDWO/2hO0x6Dm+fWdnBjWt/YmqMQcQdp
oipUE7GeOT168YrD/92F/JmEpQ/3p+3NRmh6aKt85/557NCZnRIZ7QI1b/kWv1P2EpAg6O0g/z02
nb29uXLwDyE10JL9T9J5j5Ci1pZ/4s+xVYHWZBs1mWbbxolZZM9Tx4vNqcIpANpv6hJ25fBUp0lZ
TURD9xGoTJpCEeeMxINzL03GeBG9ErHv01IDLQUyJ0zTTwiXHFTToLW/VHUVlKWZJmZPBvbErsLC
3G7TTJsgZAfl/BCCoVOWyBIWxitmHVvRrEUECFxQauIRhuC3ea9k1eF08H5r5ewiOmaeqks2Ve9k
/biOWguKJIWHZaC8NRjB4M+ncxp5fEC9z32848BAYVM6Wu5MeTtr8xpZ9tlOKSKSh3ctltN/OKfD
joxIamyMMAvGce/Hz/88SilxbM1ejANSOP8GCckxhLiqiY0FRBkMp3lJm2GN7OZ2UDtxT/hhajm9
crPCMYBVKokKRjqJgHXXb4JFW5fPc925zKleyd37Yzjo2hBQ3joYvaIb8GUmozhNbg1XvR7Ony3a
G307sf3wK4auedhfpdGtQmzdn1OWEE9AxFXXyBEIuZ254Q4mxQAvzSZ26eNygy23fLYs6xf1b8cZ
zn3k0YBE0IGYNCgl7abLvWFlY0VTfYiXvFnbseVKG4FnDwYnob/mAW+hYwnMiUMrku92xSHIKejj
3cCbgDNw94O5qQQzP9u9VfCKXliL+G9xd4W/A7DA77YyVasIOp9PygUEiw9xpxPs6RQ2F0kIUFJP
tgpcuiZWbUr5vxlv8pVhsx5NcOj+rC8xIR0y2VHKpOxpDRT+sQ3We6ykFBAvgh5cyCcPoTGRscIv
rzf2vXJmipfvKu1G5ZBGPh31FPo8jfOAWYDD+RN/gA/VW0vN3r3gyl/lZR5VJif1XtJcHfE1Ro1n
XjQjiZYJgBaXsGhp7hzRlgMhauU6xwpXoBYWxN9RfDwcODNYLb+/hyjrAuv2FyrJQveRPVFNMJ+Y
0vxom/Z3UyWuZOVfADaYKkHwkQHmVdVl+LZUkRWFk/lraFKZQQFsGV0jqaKYpejBc6aeY74I1eGZ
XdRVgvhDfKsTqvAGCK4zfOBeebkeNchnb4KNzaEQfWiGsbKcDrn7nHjpJuTd7cK0hMnSfoaSLIUJ
FLDtyOD5HGf5ZoQJZi/KBFGxhuVSWXzJ9El/tHdJtW2NUvnA7QuEPSE+O4fvkOvFVdvD8c88C5i7
/NHL9Rmg14ZurOMEVU+ACyqmvOeYdBZW+XPWlj+bMsM5lYY3IGeVi9vX//NVlesdc6N8LwztPBJH
Z0jUCnq/aUud9L4jcRJKG2w5G63xgQzHtixKwNyE/OloigJRLEehNS45jUSY25Ip8509uLO5QDKf
cdtdoqLeLcoJxxK7F1lR94q1Bys4OWz9kncmiYSIzgD9nfXYRmxNnL/swNa8G6JQ34kj6hexqELN
trlZHZH3ubKbgampQ5mH6e97V/K86n5WLrHDvnVLm3gab+7wYioxYlFAH0hIE1r9CrCZEafWN3lx
3w7rLu9JJlAHXCY1nlAuasoUCcm/DFrosPD1TDJ5aA2j8csZSeTB/Uy2biidEsmP16R1jvTddFrf
mQPrGMQolNdNYtH0tt3ETroqkt4uk37sK64d5zYzjOpmXWIKC9oVO/+q4sv9tX5uIAobHTleNzCJ
n3RUouRiPzo6T1vM/f+K3OW7h0SD2FZeJQOkA6IutaBFF8exwzyYotJiqPPz7EdEc2BNdldPNu/5
D5cWcPatfzLlGBblQlR64JdKBix49wjNn2DXsm0Qndhr/uG+vxuuK2XDwM7KUCTvrdHTW6NkRFqD
weo1hj9L7lgwGNyPtrnaWUcz4T/T8tb81Cwpfsw7Fk8QQAGgnU1jaXU5eVEuZTYJ9c6OZH6ZH1R9
u3g2GWzp98IJwsSRg8RS/w6mksqqg1KaanVqBBBmnT8U5TyDTOTkBXRIphaS5XzhMVBmxTlUcv0p
4n4iv9mKjWbrL/J8sEyYI+m609DmA9jSx1d4csuIcHfPxY8uQpVkaV657HiN+iR0eZVv9SQfM2Sx
ABH1wjX8pH7I17si0b8wTnYjJnZhkD9U1N8V3Fo2KE+L0HPXTR3ARoJXZ5vDYuc7lseoZIhG4cqi
Gy/FP8RBY6drrA6FA8og/BJfawdBFA73a1tNKMBPr06mcY3UUXTudctN/UlV8skKO9M2ADnEuvjv
jEsjmjGBnZr0zk83PRn+2BH//GVZDUVewD12QWOwYWQwWKgFZlF2IfTvY14SLCZ2Phw3DDHzZYMW
fAp7siPJR7GcwQDSGYKvrO7idWXRJaLBnhiUg14cr+W0GwkFlAp2sU5k+FHYAabzVV89jNKysrgM
knI3xZqLBIItbYxPUmUMEpCq7uCbuCevMKY21MdhzG+H7GtmdHYHe5Yu5RZpE/bYhZkYA7rvwSsW
WkF2P7vJC+FZPx0qSyoo1MV2heCRHjV+x1pHWJeM2YD1Wtuk68z1IuXo/3wCW2Ovl0L0fGzaDgl7
7gZWZwBg+jhp9ZbgT2ivtvCxLrNFg1zqjbPc1Z9XIIYC1sBxa75nVVlJ5JmHc7JgVXybB1RZ4nQA
RP4w/2/0sAZ7MGPIcZANDrUJPmY6kE1AkX/pdw4aV0xW1XcHox0GXiuPpq2tdwQ0wKqHm6z57KOS
GPedWH88avALb+5b713I+fGGIOQUidoHl8acUHWbsNuXfFNPb3TKZ1djkrU+R8WZUwvkzn+FhqSV
m86fRZpdvqvn54oAwTAzTJiuBc/CJlqSlOE+YuzJaxwoKBUZPgQH2BNh0Tf6tZwTiL1G4vriaKVK
ZqIVSis5vfyjuWb2ywl+OlK2+Mo6yU/XAo5TQ+4wXSJsmuU4UNJTqEvdslHwI6evWi/q7JA0NcMa
7qz6WI2KJP/p9fFwYn2yP7lUcNufON5UpSHsLYTrhybzst6aRYreYTkcRQ/DKqQSrF/N/Yeq6Krz
QVgFRwLfHQ+u18V8+eZHfMIPIhIctIk6jKsI9W0MOBjTEhf0iTWjBeI9+D9wtDniUTiWESK5KTad
kTkEvqko/+pnivIzqxg7N/xY2mzhGlGj1A3ZBg7Du0sA5wrVx8MWQjeaeN3ipQ7X11eyPFp4FJIz
uS7ztOwdJbWnc55fzbKV9jU5pH3RDf7qgFjj6EJciIHdFWapOsFxRemMvTeJDe2utuHBJrb/5fa1
VC+QbfIE23vOk9fTmZq/Pe8PeLJ8gZ95H6ICuH//kEDkLd98aoofa8rQP2FMACgr2Rs4mZ0zd9AI
HtVL3ZKGck3HpSum0biTHc2l7Hy+NICpa92LaTeFIhqoWuDwUotUHw5hUETtejB1qaWZHZc1NxJL
pE6oFAMliYpkg4z2HIbbGye+NZ4Yoa25SO9lVBNhBw5va+qwuBOfAJD7aUEwTTntiGUUR4S04dWf
DXzm1vSbxNx2TguZrDfApwHvMtA8nv7Bo7uINawuDTOmevDSbp8tdJg7EokPjWN1Uxa/OHXlldnD
s8dPrMy468TzTd1AS93a1vMPO6xCsGt/0bZlZib8OTgXBQb9lk45HCBcBlZrQfmpMCqLbAfi+qKc
59NVOckQc/V5ru771JwOPmDOT4Lhr94ST80iJ/AMqgDXpC4g9w+vs1FAZ3pzpwXshRcGghIjA7jU
b8XpLhaQd/PISlIEvt/pf78GKa4OzUE52dK21SfRSKe7tQAQ0oeekyR13RcnzkM2fxo4aHv+fZ4I
3lECsw/I+st8j4OsCczfK5CyjfdoiUyhhpZCYEVoP00BfiF6NeVOaj1Ol5WndKi1j6Jtz2mcWc9W
yXG7QXpcvy34cgkctjSA/l8xVGdzxcCNrOBk0zGz7XjTkn/cykjhoW+7S81nxhALHqROyYQLgXtJ
6SN+On+Da7S+Kk/R+C4hLVNnD92zKTye5jYFogJmJFB9N8Vs6coiGG6GAk3xbkSwooSc9Wc2klZG
16H6Fh1+QHDXSFSSJbVEW14QDOg4rguMIghAo/5Jo9UhriibwlPpZIkvVk21vjWJD0nbea17fy+Y
TegLKKectWdjfuhJ5+WQntSv/bWsaOQsEa9ouH0SOKnfXpkbR2r/ZkHzrraKLIWwmVs54zkX/i5d
XvdefCyj4hftTNc1fLbvdCm/7fxHbwI+f3i75T2GSPLB5HnQL1jgbBCiFe2knOmpKLBE5zOfdCDr
alFaeYLrDD8YMWyQKu5LsThzk70bEHqEDXMgERTnMrOdaTubLfFeetaLHhsrFYpBTPZdQY6eglwp
SGONLzDdNpfr/9NTXUrOxRP/B+KrVVwbBvCKVo1pt3Fmk9NCQgCd+L+tqKupSYez8l3+AgR6Bsu5
KuYnmq7DgPUrCo74eYXDptUGvJ8pcVhGnCnjauKq1qTamaL9Ga0+rO9qNcm5a3JX/D2xr2sP/xrn
RkbcKpQQphhXS9xZo2InAGbVLV5aXbHKxdaach0RxQIIvA0gHMAqcOdRmAoxsfar7c6I0r7WbVs5
dYkmxrZ/MpWobvDfoBQH4ilPaPZmZNByLTQcQWgZ1o/O4GAnaYNSfwIQ1ZWJggmptcb3f8cJjrDn
yt8J73CB8b+J6+U59EQHrf/MZEImIi3gSzsyFl3rb8enp2tE4uobVTkbAm4Y4V30AE/q8NW+cOBs
2ZZqljbES3aK1YNrHeU+34PmnkhQ1Bv96o8YKMzuaWmwNtOm3Xw3aHB5btFJCL6O0IJ3RwQt/9wE
V8Eu3WvPAVcMj9YjLk1KubD+HvVfD/AbsvC4f4eT0JcRea18CdxFnoumNSd5cgF8PYOR/+ZtUhmz
BlcwO+aLAlETyKJvVaUsaH+uFaGDhTTUP0hTmu5UOInNuI+YWwkb+DGIk5VlIqzTzMVuk4GeadVH
hBbI1Kx+ISVnVEF/Oq2SBtxA0CjFofEQrqlcNcU+fKvzAh4jRiHtA9zQvB20+SMR/GaE1ESPba98
AbMQ6UmEz+npUQtNWvl6RJ8L/FbkbXwKMTe01H83NLFAEZIVypG2v1W8BW5LHYcJRw1IQOTSDk77
zLdzpyUudEtn5tinKbGgmIrnTbQmVZiIrxFM3LpY0ktMF5McE7eamD0G9VM7BxB0G657tb1TsyH9
8L4V2OTYstwWBQis9ecaDNygwDIcSgvpuyWo0de/sUjt9SzvhXjLJbJFh9qj2AqABEJiIAK4dl0K
9ffo0a8K0TUql7gwM+WWZeK9AafSkayyhzyhX6rBgzNydD9KAd2Y1mXxgb7BoBgNKVlNSGxTNZVi
4ipbKMkrB2t0cJMV4sKbb+jUtgnayP5HReVKMwGyjOQbxX1oR1hJonKp1n1VMdsfWGW6Ejy2by0F
Gy/U7YyliuKWTGppcwi1qpGB/Kov84OjjXJVeCvRoGnJJ1UY9lHhChtnKVn3oz9qdq54xsHabZ5P
Fb/FP353AMyndl8LMbeVHIZmsSOhuDP+wV8ID2hiFO/Ot665FLV+r3UzNryj0mYuKFYkJoHTfabe
u4bJvIfmEvT7V8CeHtJQ9tmpALUTFuh7dNTa3kiqaHu1+E9rljcFjY/X1tX4xiLTcokQEuv1AyC+
JquWYqyosTTOqyKxinLGFqJEc2iqbMcMQ3l0b678njpNQ5ekg2dHN4C+1vYwTDWt79nsZAdSm9mW
Yh+Tgr3vnaB16nV4fCNXSMjDYd9gjxh2ctVS8hkHpNAKI8o4adjlR9hczReD9TZ84cdZPTyAVmQX
0wylGn7aEkjUfJn2RPxIgpSlfP/SttNEnQb88GJ3qttoogY+2szZ62XocggNQf+fMX2trRl0YK5j
etojPNqyqcffDCS6b8f48wUraC5W7dTr5VdxzEDyftKmMeLgg7MbAU1jfCULqvW2cOHsO+YfM80V
RdajTe31b1Mo8R/3b7IwHL2y7zW3EgitQeWM5E0ugYXBJWHwntMSvm7h+677T3MFMGuQd2kKx+18
CRrV3wHLGCmvvuqKtsgSV+8i5JjMZA0tVuovcwFUElC3PpZxAfXWYUZAd5JxGSQb6lVZul+Mvs0J
2qBRmMvHmhUg+sylvlX5WIj+YizfQnlwkCU3VHZF3szC2CcAR3inbIF6feAQeBEYUTF5AW2HgW63
lNLT3IW9ppye2lASdQAYRheBqjNHGQCzgmOF0nc0oGoMXgZ3f7GZUxDVz25Y3dRigP5lxh9mDPUL
HGBFbGlYTQz/H+Ih6FaratDlQRZnq+AGKJleOOmKSt4QxjopD2J9A7vlD7VAMrJSm1b2+O4a8uZr
cGBlMya0csESt4d0Tkc2MdooOZ/gpNdOJmcYxWsFiFVppSpt64Tiw7sgogez9XezPVDXr5BlwfW1
nKguPqDjmoXqIpU5wu8I/G8eayxkxQgDIBrsNRGTkP1SWYz36crHWC3zTp0U4SvMiwdkwkdwOg7h
tyujs/daWXjin/evvoOg16nIjUCWmdBcFSUN/4LxNlwAhwEM4XvhNoNtfikasElD9uLdampy7KRe
evmRgOirZhpjOM+BWhOCoPYFjj765Sovw2kSiTtJHX+GomokwBBe5eU4QrZZTAUjnLLxIyIEZA4L
9mdRPBPasIpExbAtEh5MN2Puy3Pp6xvdRomfe2dM1OMwyzJQojIPO/YqpvwrBgXKuZ4UgeZD1qvN
Sg9xz9430yAG4GbX1ygHJan6cBYZb7ex4Nx4xrXUj+JkhtG9HL/OxAsbrm4zoHsO8PyxB3TOYByw
9Ny3dBafrc5EBCZ2WF+veNR24ujMvo2IYaqHrY361/ljARO7ODjCw/COH1RJV1dSSKI4V2sDeYe/
wP+hAbpMSm7kmNgi1cn6Os9CsxVv2ejYsoB7H3+7nlz/FbB6Dk4tz+wzOyF7Yr64apHqLIVm9BRv
0JaE5drnhKkOKvPmAaajpx6GAdfCC6gtHWlZjxY+LALNLo/rCM84yxMTqvcqdWjqL5aLUCZ75wRV
qPKKb/DWBMnNmcmuMJXYnPzUDbK6QyyRyaNjTrtzMyYdi4+QO0fwLH0ONF/N22rTC69GazQzn83x
Uu6vHyExuy++LLNCI69kj8tFGFO5VscOMfZp7PZVtU48r7KvEMkS7gkIjTHgIEydGC/0djWVYqXZ
smobuwj1RcqFYyjhj99AqINtQQESb956NfUJahvRkaPX1SEbmV0iK/z0DYKT4oC3TF7QVTaCQsaD
uON05ndpSPe0o3TFcLvqwZGy5ok4YM+Khy4Feos36gHNkAvpa75OTqW50jos/FB32QQBWNznuyZX
uHzveiBk4r8g3WhgG5Wwnj/DbNvl43jZb8o27WZCh1VFX4NYqCSX/kNKgbWUfqCAIt33Xgy46Unw
mvQk/KH9j7YgaZPcbJyJDue3Ep6wXTA5Pz8TH74WSqOcZdB4E+9Coo0fjP/tpnqnb1IJvZUkUtog
VWRISU2CyaWi/4BzXWEQHZe0KVLDnisa9BT5O39yhf2BdCWS2K8e0as1W1SqgpmJ4PeNpaO+08mW
OtCs1G4Qid5F8xMgq9g+wJxzWyWETE/HQrrJj7jLX38CQwdAbaZCAEFuO1Zo0/U36kEST88uNPrL
/07lFSQP+RXq6Dm5jvjXW8A0QvuBA3WDcD0txT5URwLPt1k2SG87CWYf1kANDmArBZTS7LgksqQE
ZDDsItMHL61LnE+2Jii2uSV2x3PD7auKWKRADOXHoXdhMobMkYaqifKJa6dqSHc0IULRWgSadfJK
Ej8NkxnNhnkoql3WgHmot26ieQoHOtcOds30z8B4+zRNoObSumocqCebBlhKQMg5q6b0jYTTn+aC
vB2B4FXE2FlYLp1G/29muKaL3LTLrws5CDOg8sV7DjeVE6rBMX3W6dmLXG+7xrsHMTJCJVEuusHi
tRTNfmBB2eFLNQssHcvxvMcDaODZ3jGLjkmbEYuXA/mBiaVPgjQNdv4Uiv/tjPEXxhGsw1R1FDnf
ipK423iNjrdTg7yZQGpMCuV/A+lvqU1h0tXsL5H9S/cg7SeXPeBMgcCLwrBfq6uPRtrqMxmh0X/q
TR1gu8SlfksJ//qSuPNswC3ukD0q6DUx4cyBZrPmjJpY8ISIev9ueHMjfu5A/a7GkQdKtZ6Bmv+d
4w1OxoTsaWv4OPCp8BvPA8+lGs/qKRiKBChuhV5JEbYA6h/MMRVisbf00tBF806M9cyuY2A5Wmy6
ZU/+Q5+LmYYzR5sAjPbGzwq78YZEfkR24x27icdHNFvSCBKnAOGliqJPqDa2UIhtGymjZwoPCKoJ
yky0B4k8UaNoZO4vydJ/wBdq7YxwpU7l6f1WLTCan8xscfLpqYpj9DZowQKB6Zuy3hfp3ABQoADK
vUc7rYhetLhS0lwYrnFNH0wSrJRNCnSXTBOlhltx+E6+ySMXupkmSGzpFQmKnGB593FDGNXb02+I
fm+3DubR6iE41lOFuyxBnaNZ1zqYLC0N/kkJa9nlrIF/BIpR52pyiEv/dixyHCAHDgN31hkmoK81
HEnx6WwJBEeVmkyooweLExT+knZNwrZoE5oErgkIwDwMS1LfEVxpA8grrnFAq6fpbaPfmX/crOoQ
4F2N70TB6d8G2719Y3mypi9RC4ajIE8pbbQHqUNfmw3DJ9hyCW1xtzY1BDzH42ttPj1WRO3EUawe
o8bMVGrRPrhqOBs3ooEHHItdGJnizMKVX9MVUtTMeY+Jaer2lwf4KyzdDenDOgefxAAtIUL6Wf4G
IDtyfCcsLFm5QF1ZDEBR69ROmD8CkDQnN/hE94GFiB5CZf56rDNGou3EgtSS5Qy7HvSQiAN4WaxU
af4hnaS/1I+CNjXPgjMi09X1EXroGKfqeyK4PRGT+mxSv9ZatiOlHNJmFhgVnRXlzeqKCezt3Hxu
QPTK+nF/UqYMqUyEbfcjaIB06oqX+NZEYP4GjXDQ54n5GvlWc4kqUKApx+M1vPBpbvfxuWrMdRnd
j9ZMILJO6Qhc63RkNgCuUEY5tp84gYOH0JDGHNxtjFwv5m7RH4DOIa2KRwR+8A71C76zLPuT9/IH
6r/Z5BeVup1DY2ZGMaQtc3m5QBYiz7XiHLycChDmIm4I2UYHLtan/0MEKWcWUtske+rIHcB5e+27
cRLnMZjMaPVTpP37+jAoMU4My9/EDctyDMTxB6qU7ILNMXwsXzouP2x55CcU5bQubmIyvbNBgaZG
NnapPK/P3J8M/B2r0Xhbey03p4bN1OrM6JowayHyDYXgVzSAaXk9bXBpElqPIMO4ezc4BUxHRXIx
+jogNfrQdWjNhGKU1U9/LCgykbRs6TnMsHMqLJ6wMWnTk0nQb0dhrMftY/6Kx1nuKpzJbYM7fSDb
eJ1Pd7RHNTCYyYLv68P1lvqOGa3rVVFqgsgjeMFJs4w8rlz39wFdP8oTiOU1zcjUPl/l73BdOFzh
C26iipJfecODu8tV5pmrrlT/QtIKNhFmk2FU0Sy4lofTUZvcaZLapnAFANq6FPX4Ev9l/ChJH6ds
8ztkshc8CrIdur8xpNMj05A9XeoaGp3BNq/asRxq68O3uZ5tnqldrgW2eHLkWAlaADPPWPFETDGT
pTG0F28Pg1EE6MN2Mlyn6MeUq5xzfgGC1wmSU0sxRZQnPqC1g8MmWsOvG72xxXz8mhgUP8HONTq8
2OebY6qyRPuhP+326ZPa9l4EVcA9l8lDDATVmBCJZwWPO82tv3i3lEFczimZybO9EXqbHnBCQDi4
nHcWID8qj9NSjThj1Sr/lBUn0EDNh3nF7c9eM/3zBjKBcQ8yl+JfxP9yMwVZGLzhKn7CuoKa/GiU
BmN2lKg3+3OzNCU8YJbwuD/0Q92v7T/Y+BH1k/7aUJ0I4OmtjxPx1QQdCoTGJU70CJAvOJ2FuIc0
y9QpV3pubmo8Hg+2UxTFj+0JiLbI4cuUD0ISeANa/f9LJus1hJLimf1pLy+ew+RV1I2pSXXrDZ7L
9AKPQk1er97Sfg2dRISYtxUNQQb8KlpO2XO5wEurAg/Z9wPjbu6+JJ+k5RTu1Hsunz9vMmZclh5u
8hhtT4H72O19YToJTuYNPx4rFjspGedQJ3wiYwNWeItsk8PMe/mVzAkXdIs7LxNRBb+WEVHtlthV
JAAq7NIVfl98a2u9JupHB6aiW01pgOV7yXURLG8rnvueYzyyrD5w9NWy4SAvGU89QFYKZi/HjbkM
5E9V9jMi+lSxpLAHW/2ztNboZchGAtfkJ86x06qDx1LzAZQ3WM+qZ3leZGarmpU61w8po7bGhSHn
y+r9CTq0nXs17Z5qBYGr/tos41KcVRq0rDP7GjY/hGJq3+ziaPLAEGxdN7yXIzccg5uQPY6E5w/Z
VTXBBtkfwXfgcEiyXl8WhyUpoTgBcRs3jhCasUzXMWhIePI4m/8/enR+ut8CwEp3niTldRyGqntt
Q9h8xWPAifQVBN/6rEXyT9fG+zy/yKeV2oKj4wlIb352qEXAeAA0nzv7Sx6E2AblRKLdIcu3CpQd
prAld8vTNQ5jwfV3HuoR4q3W32Dr6ew2+NvaWht01VrS0mzhERL3J5oCyyQ0pvSk0VT6kF7AlCeI
qmZQf8DtHn/EbdDptlhTukHNot5oU3oppFn7m+JZAptMjG4KwrIyuTPOD2dvGpBU/pCHEhUV21CK
4MEGZqflwT5DyEa0cVmDsjoLniPapKB2Rvd6RsDU9K8jR9UPKAEmmebG+RZpDkuFp5q4xZPYuUPr
9R+Vifmt52LfPoM2K7x17K7jxLxnmvtvOvOTFOM2d88XaXnNYa0flhUQn+WUT4w6Rmn7UpbM+i6b
/xE6KFYB6/4WWbBe09fSaaa5p02qJtXF3zRvpvBX7LkcbkSOpbarv2CylBXxI0Hca0GvROkD1DHP
ekHFk6QBmTt9JpLn7Ixk4qjBfEJ//t+h+Mnfuc69jPvDEBdZxXEHbrWZV2WzJ8V2YzIzIjEAGgPD
gsmF0JBluTznTo+WYTvXQ8t6iEvgkbvUXRDKHFW5Mo1wcHJOhRGbf+lprbvYr04+8Jw7zVjY5pik
xXETeEnwhmCda0lkU2mYkuXRcRNYCrThb/AmJpAtFU7aH0FvoU64JI/yJ8CTyGii3Mnq5DNnGOaG
ExDYriywQZT2TPm4jeY5JHe7cQNtzivkitI/z+Bq6NM+VrkN4O393ighNwPkxE2aFr4jOBKS2A6+
bBu7YAIpo1Us3kreZUYNVGw4F6mOtfts3CZlk6pBZZZhVFY9vGyZUSURVN4rM/mZMufX4LwS+fFu
KL6AWbj5cjVWdkvWhScWIjw8qXvyx/MN7kKXFb96oKZAZnCYv3epkDyuxhPypPOFs2vKx4BkosuY
aREO0RKtCJeAyGsk3SMbbs+AUQHxCqtSJSJz7wYCvBjinJPHq63jo/KJyyRP2952L754ijbTHXrM
j0n3oT73c2DU4MaGrD1EzmiAdsDuU/ibBaVddrwoFcp698xBVBNWeALytFILztMadyQxvzQCrkKL
ZYYiEC2PF0SYUIJN9IP66fU5QompEl1Teo8ddtYeJWuZ0AGFrhSR0E+0U4nyK8F+Odhj2LQoFZuW
w40khmczuDTjSUX7Ub63TQzruYq5AvvLOFdre5fNcaEGjVLxGWnHkKk+AVkK0HtoFFAEgzBKjXv1
SVCuQ8UrmO8e7I8udNaZtTtzek1/OGrwRvqvdccc25DsqpKK0u5t4nGo+dwbAlx41aU/uMX2jxNk
7313BFyIN6W46H+EKoIOX9oKKYYSWEebQQQQBX/rFt+cv8d5mS0AFnkZ5EUzJquBTmvTKVMHWIUh
wqFaJbU5bzh6+/N8
`protect end_protected
